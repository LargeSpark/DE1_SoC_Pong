// Top.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module Top (
		input  wire        audio_refclk_clk,                //     audio_refclk.clk
		input  wire [3:0]  buttons_export,                  //          buttons.export
		inout  wire [35:0] gpio0_export,                    //            gpio0.export
		inout  wire [35:0] gpio1_export,                    //            gpio1.export
		output wire [6:0]  hex0_export,                     //             hex0.export
		output wire [6:0]  hex1_export,                     //             hex1.export
		output wire [6:0]  hex2_export,                     //             hex2.export
		output wire [6:0]  hex3_export,                     //             hex3.export
		output wire [6:0]  hex4_export,                     //             hex4.export
		output wire [6:0]  hex5_export,                     //             hex5.export
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //           hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //                 .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //                 .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //                 .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //                 .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //                 .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //                 .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //                 .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //                 .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //                 .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //                 .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //                 .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //                 .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //                 .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //                 .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //                 .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //                 .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //                 .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //                 .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //                 .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //                 .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //                 .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //                 .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //                 .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //                 .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //                 .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //                 .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //                 .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //                 .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //                 .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //                 .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //                 .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //                 .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //                 .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //                 .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //                 .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //                 .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //                 .hps_io_usb1_inst_NXT
		output wire        hps_io_hps_io_spim1_inst_CLK,    //                 .hps_io_spim1_inst_CLK
		output wire        hps_io_hps_io_spim1_inst_MOSI,   //                 .hps_io_spim1_inst_MOSI
		input  wire        hps_io_hps_io_spim1_inst_MISO,   //                 .hps_io_spim1_inst_MISO
		output wire        hps_io_hps_io_spim1_inst_SS0,    //                 .hps_io_spim1_inst_SS0
		input  wire        hps_io_hps_io_uart0_inst_RX,     //                 .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //                 .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //                 .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //                 .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //                 .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //                 .hps_io_i2c1_inst_SCL
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //                 .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,  //                 .hps_io_gpio_inst_GPIO35
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //                 .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //                 .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //                 .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO53,  //                 .hps_io_gpio_inst_GPIO53
		inout  wire        hps_io_hps_io_gpio_inst_GPIO54,  //                 .hps_io_gpio_inst_GPIO54
		inout  wire        hps_io_hps_io_gpio_inst_GPIO61,  //                 .hps_io_gpio_inst_GPIO61
		output wire        irda_uart_tx,                    //        irda_uart.tx
		input  wire        irda_uart_rx,                    //                 .rx
		output wire [9:0]  leds_export,                     //             leds.export
		output wire [14:0] memory_mem_a,                    //           memory.mem_a
		output wire [2:0]  memory_mem_ba,                   //                 .mem_ba
		output wire        memory_mem_ck,                   //                 .mem_ck
		output wire        memory_mem_ck_n,                 //                 .mem_ck_n
		output wire        memory_mem_cke,                  //                 .mem_cke
		output wire        memory_mem_cs_n,                 //                 .mem_cs_n
		output wire        memory_mem_ras_n,                //                 .mem_ras_n
		output wire        memory_mem_cas_n,                //                 .mem_cas_n
		output wire        memory_mem_we_n,                 //                 .mem_we_n
		output wire        memory_mem_reset_n,              //                 .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                   //                 .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                  //                 .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                //                 .mem_dqs_n
		output wire        memory_mem_odt,                  //                 .mem_odt
		output wire [3:0]  memory_mem_dm,                   //                 .mem_dm
		input  wire        memory_oct_rzqin,                //                 .oct_rzqin
		inout  wire        ps2_0_CLK,                       //            ps2_0.CLK
		inout  wire        ps2_0_DAT,                       //                 .DAT
		inout  wire        ps2_1_CLK,                       //            ps2_1.CLK
		inout  wire        ps2_1_DAT,                       //                 .DAT
		output wire [12:0] sdram_addr,                      //            sdram.addr
		output wire [1:0]  sdram_ba,                        //                 .ba
		output wire        sdram_cas_n,                     //                 .cas_n
		output wire        sdram_cke,                       //                 .cke
		output wire        sdram_cs_n,                      //                 .cs_n
		inout  wire [15:0] sdram_dq,                        //                 .dq
		output wire [1:0]  sdram_dqm,                       //                 .dqm
		output wire        sdram_ras_n,                     //                 .ras_n
		output wire        sdram_we_n,                      //                 .we_n
		output wire        sdram_clk_clk,                   //        sdram_clk.clk
		input  wire [9:0]  switches_export,                 //         switches.export
		input  wire        system_ref_clk_clk,              //   system_ref_clk.clk
		input  wire        system_ref_reset_reset,          // system_ref_reset.reset
		output wire        vga_CLK,                         //              vga.CLK
		output wire        vga_HS,                          //                 .HS
		output wire        vga_VS,                          //                 .VS
		output wire        vga_BLANK,                       //                 .BLANK
		output wire        vga_SYNC,                        //                 .SYNC
		output wire [7:0]  vga_R,                           //                 .R
		output wire [7:0]  vga_G,                           //                 .G
		output wire [7:0]  vga_B,                           //                 .B
		input  wire        vga_refclk_clk,                  //       vga_refclk.clk
		input  wire        wm8731_bclk,                     //           wm8731.bclk
		input  wire        wm8731_adclrck,                  //                 .adclrck
		input  wire        wm8731_adcdat,                   //                 .adcdat
		input  wire        wm8731_daclrck,                  //                 .daclrck
		output wire        wm8731_dacdat,                   //                 .dacdat
		output wire        wm8731_xck_clk                   //       wm8731_xck.clk
	);

	wire          ioperipherals_ddr_read_waitrequest;                                  // arm_hps:f2h_sdram0_WAITREQUEST -> IOPeripherals:ddr_read_waitrequest
	wire  [127:0] ioperipherals_ddr_read_readdata;                                     // arm_hps:f2h_sdram0_READDATA -> IOPeripherals:ddr_read_readdata
	wire          ioperipherals_ddr_read_read;                                         // IOPeripherals:ddr_read_read -> arm_hps:f2h_sdram0_READ
	wire   [27:0] ioperipherals_ddr_read_address;                                      // IOPeripherals:ddr_read_address -> arm_hps:f2h_sdram0_ADDRESS
	wire          ioperipherals_ddr_read_readdatavalid;                                // arm_hps:f2h_sdram0_READDATAVALID -> IOPeripherals:ddr_read_readdatavalid
	wire    [7:0] ioperipherals_ddr_read_burstcount;                                   // IOPeripherals:ddr_read_burstcount -> arm_hps:f2h_sdram0_BURSTCOUNT
	wire          ioperipherals_ddr_write_waitrequest;                                 // arm_hps:f2h_sdram1_WAITREQUEST -> IOPeripherals:ddr_write_waitrequest
	wire   [15:0] ioperipherals_ddr_write_byteenable;                                  // IOPeripherals:ddr_write_byteenable -> arm_hps:f2h_sdram1_BYTEENABLE
	wire   [27:0] ioperipherals_ddr_write_address;                                     // IOPeripherals:ddr_write_address -> arm_hps:f2h_sdram1_ADDRESS
	wire          ioperipherals_ddr_write_write;                                       // IOPeripherals:ddr_write_write -> arm_hps:f2h_sdram1_WRITE
	wire  [127:0] ioperipherals_ddr_write_writedata;                                   // IOPeripherals:ddr_write_writedata -> arm_hps:f2h_sdram1_WRITEDATA
	wire    [7:0] ioperipherals_ddr_write_burstcount;                                  // IOPeripherals:ddr_write_burstcount -> arm_hps:f2h_sdram1_BURSTCOUNT
	wire          system_ref_pll_outclk0_clk;                                          // system_ref_pll:outclk_0 -> [AudioSubsystem:clk_clk, IOPeripherals:sys_clk_clk, VGASubsystem:sys_clk_clk, arm_hps:f2h_axi_clk, arm_hps:f2h_sdram0_clk, arm_hps:f2h_sdram1_clk, arm_hps:h2f_axi_clk, arm_hps:h2f_lw_axi_clk, baremetal:clk, interval_timer:clk, jtag_fpga:clk_clk, jtag_hps:clk_clk, mm_interconnect_2:system_ref_pll_outclk0_clk, mm_interconnect_3:system_ref_pll_outclk0_clk, ocram:clk, rst_controller:clk, rst_controller_001:clk, sdram:clk, sysid:clock, system_reset:clk]
	wire          boot_from_fpga_constant_boot_from_fpga_on_failure;                   // boot_from_fpga:boot_from_fpga_on_failure -> arm_hps:f2h_boot_from_fpga_on_failure
	wire          boot_from_fpga_constant_boot_from_fpga_ready;                        // boot_from_fpga:boot_from_fpga_ready -> arm_hps:f2h_boot_from_fpga_ready
	wire          system_ref_pll_locked_export;                                        // system_ref_pll:locked -> pll_locked:locked
	wire          arm_hps_h2f_reset_reset;                                             // arm_hps:h2f_rst_n -> [rst_controller_001:reset_in0, system_reset:reset_in1]
	wire          pll_locked_reset_reset;                                              // pll_locked:reset_n -> system_reset:reset_in0
	wire          system_reset_reset_out_reset;                                        // system_reset:reset_out -> [VGASubsystem:sys_reset_reset_n, VGASubsystem:vga_pll_ref_reset_reset, jtag_fpga:clk_reset_reset, jtag_hps:clk_reset_reset, rst_controller:reset_in0]
	wire    [1:0] arm_hps_h2f_axi_master_awburst;                                      // arm_hps:h2f_AWBURST -> mm_interconnect_2:arm_hps_h2f_axi_master_awburst
	wire    [3:0] arm_hps_h2f_axi_master_arlen;                                        // arm_hps:h2f_ARLEN -> mm_interconnect_2:arm_hps_h2f_axi_master_arlen
	wire   [15:0] arm_hps_h2f_axi_master_wstrb;                                        // arm_hps:h2f_WSTRB -> mm_interconnect_2:arm_hps_h2f_axi_master_wstrb
	wire          arm_hps_h2f_axi_master_wready;                                       // mm_interconnect_2:arm_hps_h2f_axi_master_wready -> arm_hps:h2f_WREADY
	wire   [11:0] arm_hps_h2f_axi_master_rid;                                          // mm_interconnect_2:arm_hps_h2f_axi_master_rid -> arm_hps:h2f_RID
	wire          arm_hps_h2f_axi_master_rready;                                       // arm_hps:h2f_RREADY -> mm_interconnect_2:arm_hps_h2f_axi_master_rready
	wire    [3:0] arm_hps_h2f_axi_master_awlen;                                        // arm_hps:h2f_AWLEN -> mm_interconnect_2:arm_hps_h2f_axi_master_awlen
	wire   [11:0] arm_hps_h2f_axi_master_wid;                                          // arm_hps:h2f_WID -> mm_interconnect_2:arm_hps_h2f_axi_master_wid
	wire    [3:0] arm_hps_h2f_axi_master_arcache;                                      // arm_hps:h2f_ARCACHE -> mm_interconnect_2:arm_hps_h2f_axi_master_arcache
	wire          arm_hps_h2f_axi_master_wvalid;                                       // arm_hps:h2f_WVALID -> mm_interconnect_2:arm_hps_h2f_axi_master_wvalid
	wire   [29:0] arm_hps_h2f_axi_master_araddr;                                       // arm_hps:h2f_ARADDR -> mm_interconnect_2:arm_hps_h2f_axi_master_araddr
	wire    [2:0] arm_hps_h2f_axi_master_arprot;                                       // arm_hps:h2f_ARPROT -> mm_interconnect_2:arm_hps_h2f_axi_master_arprot
	wire    [2:0] arm_hps_h2f_axi_master_awprot;                                       // arm_hps:h2f_AWPROT -> mm_interconnect_2:arm_hps_h2f_axi_master_awprot
	wire  [127:0] arm_hps_h2f_axi_master_wdata;                                        // arm_hps:h2f_WDATA -> mm_interconnect_2:arm_hps_h2f_axi_master_wdata
	wire          arm_hps_h2f_axi_master_arvalid;                                      // arm_hps:h2f_ARVALID -> mm_interconnect_2:arm_hps_h2f_axi_master_arvalid
	wire    [3:0] arm_hps_h2f_axi_master_awcache;                                      // arm_hps:h2f_AWCACHE -> mm_interconnect_2:arm_hps_h2f_axi_master_awcache
	wire   [11:0] arm_hps_h2f_axi_master_arid;                                         // arm_hps:h2f_ARID -> mm_interconnect_2:arm_hps_h2f_axi_master_arid
	wire    [1:0] arm_hps_h2f_axi_master_arlock;                                       // arm_hps:h2f_ARLOCK -> mm_interconnect_2:arm_hps_h2f_axi_master_arlock
	wire    [1:0] arm_hps_h2f_axi_master_awlock;                                       // arm_hps:h2f_AWLOCK -> mm_interconnect_2:arm_hps_h2f_axi_master_awlock
	wire   [29:0] arm_hps_h2f_axi_master_awaddr;                                       // arm_hps:h2f_AWADDR -> mm_interconnect_2:arm_hps_h2f_axi_master_awaddr
	wire    [1:0] arm_hps_h2f_axi_master_bresp;                                        // mm_interconnect_2:arm_hps_h2f_axi_master_bresp -> arm_hps:h2f_BRESP
	wire          arm_hps_h2f_axi_master_arready;                                      // mm_interconnect_2:arm_hps_h2f_axi_master_arready -> arm_hps:h2f_ARREADY
	wire  [127:0] arm_hps_h2f_axi_master_rdata;                                        // mm_interconnect_2:arm_hps_h2f_axi_master_rdata -> arm_hps:h2f_RDATA
	wire          arm_hps_h2f_axi_master_awready;                                      // mm_interconnect_2:arm_hps_h2f_axi_master_awready -> arm_hps:h2f_AWREADY
	wire    [1:0] arm_hps_h2f_axi_master_arburst;                                      // arm_hps:h2f_ARBURST -> mm_interconnect_2:arm_hps_h2f_axi_master_arburst
	wire    [2:0] arm_hps_h2f_axi_master_arsize;                                       // arm_hps:h2f_ARSIZE -> mm_interconnect_2:arm_hps_h2f_axi_master_arsize
	wire          arm_hps_h2f_axi_master_bready;                                       // arm_hps:h2f_BREADY -> mm_interconnect_2:arm_hps_h2f_axi_master_bready
	wire          arm_hps_h2f_axi_master_rlast;                                        // mm_interconnect_2:arm_hps_h2f_axi_master_rlast -> arm_hps:h2f_RLAST
	wire          arm_hps_h2f_axi_master_wlast;                                        // arm_hps:h2f_WLAST -> mm_interconnect_2:arm_hps_h2f_axi_master_wlast
	wire    [1:0] arm_hps_h2f_axi_master_rresp;                                        // mm_interconnect_2:arm_hps_h2f_axi_master_rresp -> arm_hps:h2f_RRESP
	wire   [11:0] arm_hps_h2f_axi_master_awid;                                         // arm_hps:h2f_AWID -> mm_interconnect_2:arm_hps_h2f_axi_master_awid
	wire   [11:0] arm_hps_h2f_axi_master_bid;                                          // mm_interconnect_2:arm_hps_h2f_axi_master_bid -> arm_hps:h2f_BID
	wire          arm_hps_h2f_axi_master_bvalid;                                       // mm_interconnect_2:arm_hps_h2f_axi_master_bvalid -> arm_hps:h2f_BVALID
	wire    [2:0] arm_hps_h2f_axi_master_awsize;                                       // arm_hps:h2f_AWSIZE -> mm_interconnect_2:arm_hps_h2f_axi_master_awsize
	wire          arm_hps_h2f_axi_master_awvalid;                                      // arm_hps:h2f_AWVALID -> mm_interconnect_2:arm_hps_h2f_axi_master_awvalid
	wire          arm_hps_h2f_axi_master_rvalid;                                       // mm_interconnect_2:arm_hps_h2f_axi_master_rvalid -> arm_hps:h2f_RVALID
	wire   [31:0] jtag_fpga_master_readdata;                                           // mm_interconnect_2:jtag_fpga_master_readdata -> jtag_fpga:master_readdata
	wire          jtag_fpga_master_waitrequest;                                        // mm_interconnect_2:jtag_fpga_master_waitrequest -> jtag_fpga:master_waitrequest
	wire   [31:0] jtag_fpga_master_address;                                            // jtag_fpga:master_address -> mm_interconnect_2:jtag_fpga_master_address
	wire          jtag_fpga_master_read;                                               // jtag_fpga:master_read -> mm_interconnect_2:jtag_fpga_master_read
	wire    [3:0] jtag_fpga_master_byteenable;                                         // jtag_fpga:master_byteenable -> mm_interconnect_2:jtag_fpga_master_byteenable
	wire          jtag_fpga_master_readdatavalid;                                      // mm_interconnect_2:jtag_fpga_master_readdatavalid -> jtag_fpga:master_readdatavalid
	wire          jtag_fpga_master_write;                                              // jtag_fpga:master_write -> mm_interconnect_2:jtag_fpga_master_write
	wire   [31:0] jtag_fpga_master_writedata;                                          // jtag_fpga:master_writedata -> mm_interconnect_2:jtag_fpga_master_writedata
	wire    [1:0] arm_hps_h2f_lw_axi_master_awburst;                                   // arm_hps:h2f_lw_AWBURST -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awburst
	wire    [3:0] arm_hps_h2f_lw_axi_master_arlen;                                     // arm_hps:h2f_lw_ARLEN -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arlen
	wire    [3:0] arm_hps_h2f_lw_axi_master_wstrb;                                     // arm_hps:h2f_lw_WSTRB -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_wstrb
	wire          arm_hps_h2f_lw_axi_master_wready;                                    // mm_interconnect_2:arm_hps_h2f_lw_axi_master_wready -> arm_hps:h2f_lw_WREADY
	wire   [11:0] arm_hps_h2f_lw_axi_master_rid;                                       // mm_interconnect_2:arm_hps_h2f_lw_axi_master_rid -> arm_hps:h2f_lw_RID
	wire          arm_hps_h2f_lw_axi_master_rready;                                    // arm_hps:h2f_lw_RREADY -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_rready
	wire    [3:0] arm_hps_h2f_lw_axi_master_awlen;                                     // arm_hps:h2f_lw_AWLEN -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awlen
	wire   [11:0] arm_hps_h2f_lw_axi_master_wid;                                       // arm_hps:h2f_lw_WID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_wid
	wire    [3:0] arm_hps_h2f_lw_axi_master_arcache;                                   // arm_hps:h2f_lw_ARCACHE -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arcache
	wire          arm_hps_h2f_lw_axi_master_wvalid;                                    // arm_hps:h2f_lw_WVALID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_wvalid
	wire   [20:0] arm_hps_h2f_lw_axi_master_araddr;                                    // arm_hps:h2f_lw_ARADDR -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_araddr
	wire    [2:0] arm_hps_h2f_lw_axi_master_arprot;                                    // arm_hps:h2f_lw_ARPROT -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arprot
	wire    [2:0] arm_hps_h2f_lw_axi_master_awprot;                                    // arm_hps:h2f_lw_AWPROT -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awprot
	wire   [31:0] arm_hps_h2f_lw_axi_master_wdata;                                     // arm_hps:h2f_lw_WDATA -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_wdata
	wire          arm_hps_h2f_lw_axi_master_arvalid;                                   // arm_hps:h2f_lw_ARVALID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arvalid
	wire    [3:0] arm_hps_h2f_lw_axi_master_awcache;                                   // arm_hps:h2f_lw_AWCACHE -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awcache
	wire   [11:0] arm_hps_h2f_lw_axi_master_arid;                                      // arm_hps:h2f_lw_ARID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arid
	wire    [1:0] arm_hps_h2f_lw_axi_master_arlock;                                    // arm_hps:h2f_lw_ARLOCK -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arlock
	wire    [1:0] arm_hps_h2f_lw_axi_master_awlock;                                    // arm_hps:h2f_lw_AWLOCK -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awlock
	wire   [20:0] arm_hps_h2f_lw_axi_master_awaddr;                                    // arm_hps:h2f_lw_AWADDR -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awaddr
	wire    [1:0] arm_hps_h2f_lw_axi_master_bresp;                                     // mm_interconnect_2:arm_hps_h2f_lw_axi_master_bresp -> arm_hps:h2f_lw_BRESP
	wire          arm_hps_h2f_lw_axi_master_arready;                                   // mm_interconnect_2:arm_hps_h2f_lw_axi_master_arready -> arm_hps:h2f_lw_ARREADY
	wire   [31:0] arm_hps_h2f_lw_axi_master_rdata;                                     // mm_interconnect_2:arm_hps_h2f_lw_axi_master_rdata -> arm_hps:h2f_lw_RDATA
	wire          arm_hps_h2f_lw_axi_master_awready;                                   // mm_interconnect_2:arm_hps_h2f_lw_axi_master_awready -> arm_hps:h2f_lw_AWREADY
	wire    [1:0] arm_hps_h2f_lw_axi_master_arburst;                                   // arm_hps:h2f_lw_ARBURST -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arburst
	wire    [2:0] arm_hps_h2f_lw_axi_master_arsize;                                    // arm_hps:h2f_lw_ARSIZE -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_arsize
	wire          arm_hps_h2f_lw_axi_master_bready;                                    // arm_hps:h2f_lw_BREADY -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_bready
	wire          arm_hps_h2f_lw_axi_master_rlast;                                     // mm_interconnect_2:arm_hps_h2f_lw_axi_master_rlast -> arm_hps:h2f_lw_RLAST
	wire          arm_hps_h2f_lw_axi_master_wlast;                                     // arm_hps:h2f_lw_WLAST -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_wlast
	wire    [1:0] arm_hps_h2f_lw_axi_master_rresp;                                     // mm_interconnect_2:arm_hps_h2f_lw_axi_master_rresp -> arm_hps:h2f_lw_RRESP
	wire   [11:0] arm_hps_h2f_lw_axi_master_awid;                                      // arm_hps:h2f_lw_AWID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awid
	wire   [11:0] arm_hps_h2f_lw_axi_master_bid;                                       // mm_interconnect_2:arm_hps_h2f_lw_axi_master_bid -> arm_hps:h2f_lw_BID
	wire          arm_hps_h2f_lw_axi_master_bvalid;                                    // mm_interconnect_2:arm_hps_h2f_lw_axi_master_bvalid -> arm_hps:h2f_lw_BVALID
	wire    [2:0] arm_hps_h2f_lw_axi_master_awsize;                                    // arm_hps:h2f_lw_AWSIZE -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awsize
	wire          arm_hps_h2f_lw_axi_master_awvalid;                                   // arm_hps:h2f_lw_AWVALID -> mm_interconnect_2:arm_hps_h2f_lw_axi_master_awvalid
	wire          arm_hps_h2f_lw_axi_master_rvalid;                                    // mm_interconnect_2:arm_hps_h2f_lw_axi_master_rvalid -> arm_hps:h2f_lw_RVALID
	wire          vgasubsystem_pixel_dma_master_waitrequest;                           // mm_interconnect_2:VGASubsystem_pixel_dma_master_waitrequest -> VGASubsystem:pixel_dma_master_waitrequest
	wire   [15:0] vgasubsystem_pixel_dma_master_readdata;                              // mm_interconnect_2:VGASubsystem_pixel_dma_master_readdata -> VGASubsystem:pixel_dma_master_readdata
	wire   [31:0] vgasubsystem_pixel_dma_master_address;                               // VGASubsystem:pixel_dma_master_address -> mm_interconnect_2:VGASubsystem_pixel_dma_master_address
	wire          vgasubsystem_pixel_dma_master_read;                                  // VGASubsystem:pixel_dma_master_read -> mm_interconnect_2:VGASubsystem_pixel_dma_master_read
	wire          vgasubsystem_pixel_dma_master_readdatavalid;                         // mm_interconnect_2:VGASubsystem_pixel_dma_master_readdatavalid -> VGASubsystem:pixel_dma_master_readdatavalid
	wire          vgasubsystem_pixel_dma_master_lock;                                  // VGASubsystem:pixel_dma_master_lock -> mm_interconnect_2:VGASubsystem_pixel_dma_master_lock
	wire          mm_interconnect_2_vgasubsystem_char_buffer_slave_chipselect;         // mm_interconnect_2:VGASubsystem_char_buffer_slave_chipselect -> VGASubsystem:char_buffer_slave_chipselect
	wire    [7:0] mm_interconnect_2_vgasubsystem_char_buffer_slave_readdata;           // VGASubsystem:char_buffer_slave_readdata -> mm_interconnect_2:VGASubsystem_char_buffer_slave_readdata
	wire          mm_interconnect_2_vgasubsystem_char_buffer_slave_waitrequest;        // VGASubsystem:char_buffer_slave_waitrequest -> mm_interconnect_2:VGASubsystem_char_buffer_slave_waitrequest
	wire   [12:0] mm_interconnect_2_vgasubsystem_char_buffer_slave_address;            // mm_interconnect_2:VGASubsystem_char_buffer_slave_address -> VGASubsystem:char_buffer_slave_address
	wire          mm_interconnect_2_vgasubsystem_char_buffer_slave_read;               // mm_interconnect_2:VGASubsystem_char_buffer_slave_read -> VGASubsystem:char_buffer_slave_read
	wire    [0:0] mm_interconnect_2_vgasubsystem_char_buffer_slave_byteenable;         // mm_interconnect_2:VGASubsystem_char_buffer_slave_byteenable -> VGASubsystem:char_buffer_slave_byteenable
	wire          mm_interconnect_2_vgasubsystem_char_buffer_slave_write;              // mm_interconnect_2:VGASubsystem_char_buffer_slave_write -> VGASubsystem:char_buffer_slave_write
	wire    [7:0] mm_interconnect_2_vgasubsystem_char_buffer_slave_writedata;          // mm_interconnect_2:VGASubsystem_char_buffer_slave_writedata -> VGASubsystem:char_buffer_slave_writedata
	wire          mm_interconnect_2_ocram_s1_chipselect;                               // mm_interconnect_2:ocram_s1_chipselect -> ocram:chipselect
	wire   [31:0] mm_interconnect_2_ocram_s1_readdata;                                 // ocram:readdata -> mm_interconnect_2:ocram_s1_readdata
	wire   [11:0] mm_interconnect_2_ocram_s1_address;                                  // mm_interconnect_2:ocram_s1_address -> ocram:address
	wire    [3:0] mm_interconnect_2_ocram_s1_byteenable;                               // mm_interconnect_2:ocram_s1_byteenable -> ocram:byteenable
	wire          mm_interconnect_2_ocram_s1_write;                                    // mm_interconnect_2:ocram_s1_write -> ocram:write
	wire   [31:0] mm_interconnect_2_ocram_s1_writedata;                                // mm_interconnect_2:ocram_s1_writedata -> ocram:writedata
	wire          mm_interconnect_2_ocram_s1_clken;                                    // mm_interconnect_2:ocram_s1_clken -> ocram:clken
	wire          mm_interconnect_2_sdram_s1_chipselect;                               // mm_interconnect_2:sdram_s1_chipselect -> sdram:az_cs
	wire   [15:0] mm_interconnect_2_sdram_s1_readdata;                                 // sdram:za_data -> mm_interconnect_2:sdram_s1_readdata
	wire          mm_interconnect_2_sdram_s1_waitrequest;                              // sdram:za_waitrequest -> mm_interconnect_2:sdram_s1_waitrequest
	wire   [24:0] mm_interconnect_2_sdram_s1_address;                                  // mm_interconnect_2:sdram_s1_address -> sdram:az_addr
	wire          mm_interconnect_2_sdram_s1_read;                                     // mm_interconnect_2:sdram_s1_read -> sdram:az_rd_n
	wire    [1:0] mm_interconnect_2_sdram_s1_byteenable;                               // mm_interconnect_2:sdram_s1_byteenable -> sdram:az_be_n
	wire          mm_interconnect_2_sdram_s1_readdatavalid;                            // sdram:za_valid -> mm_interconnect_2:sdram_s1_readdatavalid
	wire          mm_interconnect_2_sdram_s1_write;                                    // mm_interconnect_2:sdram_s1_write -> sdram:az_wr_n
	wire   [15:0] mm_interconnect_2_sdram_s1_writedata;                                // mm_interconnect_2:sdram_s1_writedata -> sdram:az_data
	wire          mm_interconnect_2_baremetal_s1_chipselect;                           // mm_interconnect_2:baremetal_s1_chipselect -> baremetal:chipselect
	wire   [31:0] mm_interconnect_2_baremetal_s1_readdata;                             // baremetal:readdata -> mm_interconnect_2:baremetal_s1_readdata
	wire   [13:0] mm_interconnect_2_baremetal_s1_address;                              // mm_interconnect_2:baremetal_s1_address -> baremetal:address
	wire    [3:0] mm_interconnect_2_baremetal_s1_byteenable;                           // mm_interconnect_2:baremetal_s1_byteenable -> baremetal:byteenable
	wire          mm_interconnect_2_baremetal_s1_write;                                // mm_interconnect_2:baremetal_s1_write -> baremetal:write
	wire   [31:0] mm_interconnect_2_baremetal_s1_writedata;                            // mm_interconnect_2:baremetal_s1_writedata -> baremetal:writedata
	wire          mm_interconnect_2_baremetal_s1_clken;                                // mm_interconnect_2:baremetal_s1_clken -> baremetal:clken
	wire          mm_interconnect_2_vgasubsystem_char_buffer_control_slave_chipselect; // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_chipselect -> VGASubsystem:char_buffer_control_slave_chipselect
	wire   [31:0] mm_interconnect_2_vgasubsystem_char_buffer_control_slave_readdata;   // VGASubsystem:char_buffer_control_slave_readdata -> mm_interconnect_2:VGASubsystem_char_buffer_control_slave_readdata
	wire    [0:0] mm_interconnect_2_vgasubsystem_char_buffer_control_slave_address;    // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_address -> VGASubsystem:char_buffer_control_slave_address
	wire          mm_interconnect_2_vgasubsystem_char_buffer_control_slave_read;       // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_read -> VGASubsystem:char_buffer_control_slave_read
	wire    [3:0] mm_interconnect_2_vgasubsystem_char_buffer_control_slave_byteenable; // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_byteenable -> VGASubsystem:char_buffer_control_slave_byteenable
	wire          mm_interconnect_2_vgasubsystem_char_buffer_control_slave_write;      // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_write -> VGASubsystem:char_buffer_control_slave_write
	wire   [31:0] mm_interconnect_2_vgasubsystem_char_buffer_control_slave_writedata;  // mm_interconnect_2:VGASubsystem_char_buffer_control_slave_writedata -> VGASubsystem:char_buffer_control_slave_writedata
	wire   [31:0] mm_interconnect_2_sysid_control_slave_readdata;                      // sysid:readdata -> mm_interconnect_2:sysid_control_slave_readdata
	wire    [0:0] mm_interconnect_2_sysid_control_slave_address;                       // mm_interconnect_2:sysid_control_slave_address -> sysid:address
	wire          mm_interconnect_2_audiosubsystem_csr_chipselect;                     // mm_interconnect_2:AudioSubsystem_csr_chipselect -> AudioSubsystem:csr_chipselect
	wire   [31:0] mm_interconnect_2_audiosubsystem_csr_readdata;                       // AudioSubsystem:csr_readdata -> mm_interconnect_2:AudioSubsystem_csr_readdata
	wire    [2:0] mm_interconnect_2_audiosubsystem_csr_address;                        // mm_interconnect_2:AudioSubsystem_csr_address -> AudioSubsystem:csr_address
	wire          mm_interconnect_2_audiosubsystem_csr_read;                           // mm_interconnect_2:AudioSubsystem_csr_read -> AudioSubsystem:csr_read
	wire    [3:0] mm_interconnect_2_audiosubsystem_csr_byteenable;                     // mm_interconnect_2:AudioSubsystem_csr_byteenable -> AudioSubsystem:csr_byteenable
	wire          mm_interconnect_2_audiosubsystem_csr_write;                          // mm_interconnect_2:AudioSubsystem_csr_write -> AudioSubsystem:csr_write
	wire   [31:0] mm_interconnect_2_audiosubsystem_csr_writedata;                      // mm_interconnect_2:AudioSubsystem_csr_writedata -> AudioSubsystem:csr_writedata
	wire   [31:0] mm_interconnect_2_ioperipherals_peripheral_map_readdata;             // IOPeripherals:peripheral_map_readdata -> mm_interconnect_2:IOPeripherals_peripheral_map_readdata
	wire          mm_interconnect_2_ioperipherals_peripheral_map_waitrequest;          // IOPeripherals:peripheral_map_waitrequest -> mm_interconnect_2:IOPeripherals_peripheral_map_waitrequest
	wire          mm_interconnect_2_ioperipherals_peripheral_map_debugaccess;          // mm_interconnect_2:IOPeripherals_peripheral_map_debugaccess -> IOPeripherals:peripheral_map_debugaccess
	wire   [10:0] mm_interconnect_2_ioperipherals_peripheral_map_address;              // mm_interconnect_2:IOPeripherals_peripheral_map_address -> IOPeripherals:peripheral_map_address
	wire          mm_interconnect_2_ioperipherals_peripheral_map_read;                 // mm_interconnect_2:IOPeripherals_peripheral_map_read -> IOPeripherals:peripheral_map_read
	wire    [3:0] mm_interconnect_2_ioperipherals_peripheral_map_byteenable;           // mm_interconnect_2:IOPeripherals_peripheral_map_byteenable -> IOPeripherals:peripheral_map_byteenable
	wire          mm_interconnect_2_ioperipherals_peripheral_map_readdatavalid;        // IOPeripherals:peripheral_map_readdatavalid -> mm_interconnect_2:IOPeripherals_peripheral_map_readdatavalid
	wire          mm_interconnect_2_ioperipherals_peripheral_map_write;                // mm_interconnect_2:IOPeripherals_peripheral_map_write -> IOPeripherals:peripheral_map_write
	wire   [31:0] mm_interconnect_2_ioperipherals_peripheral_map_writedata;            // mm_interconnect_2:IOPeripherals_peripheral_map_writedata -> IOPeripherals:peripheral_map_writedata
	wire    [0:0] mm_interconnect_2_ioperipherals_peripheral_map_burstcount;           // mm_interconnect_2:IOPeripherals_peripheral_map_burstcount -> IOPeripherals:peripheral_map_burstcount
	wire   [31:0] mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_readdata;     // VGASubsystem:pixel_dma_control_slave_readdata -> mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_readdata
	wire    [1:0] mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_address;      // mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_address -> VGASubsystem:pixel_dma_control_slave_address
	wire          mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_read;         // mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_read -> VGASubsystem:pixel_dma_control_slave_read
	wire    [3:0] mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_byteenable;   // mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_byteenable -> VGASubsystem:pixel_dma_control_slave_byteenable
	wire          mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_write;        // mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_write -> VGASubsystem:pixel_dma_control_slave_write
	wire   [31:0] mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_writedata;    // mm_interconnect_2:VGASubsystem_pixel_dma_control_slave_writedata -> VGASubsystem:pixel_dma_control_slave_writedata
	wire          mm_interconnect_2_interval_timer_s1_chipselect;                      // mm_interconnect_2:interval_timer_s1_chipselect -> interval_timer:chipselect
	wire   [15:0] mm_interconnect_2_interval_timer_s1_readdata;                        // interval_timer:readdata -> mm_interconnect_2:interval_timer_s1_readdata
	wire    [2:0] mm_interconnect_2_interval_timer_s1_address;                         // mm_interconnect_2:interval_timer_s1_address -> interval_timer:address
	wire          mm_interconnect_2_interval_timer_s1_write;                           // mm_interconnect_2:interval_timer_s1_write -> interval_timer:write_n
	wire   [15:0] mm_interconnect_2_interval_timer_s1_writedata;                       // mm_interconnect_2:interval_timer_s1_writedata -> interval_timer:writedata
	wire          mm_interconnect_2_ocram_s2_chipselect;                               // mm_interconnect_2:ocram_s2_chipselect -> ocram:chipselect2
	wire   [31:0] mm_interconnect_2_ocram_s2_readdata;                                 // ocram:readdata2 -> mm_interconnect_2:ocram_s2_readdata
	wire   [11:0] mm_interconnect_2_ocram_s2_address;                                  // mm_interconnect_2:ocram_s2_address -> ocram:address2
	wire    [3:0] mm_interconnect_2_ocram_s2_byteenable;                               // mm_interconnect_2:ocram_s2_byteenable -> ocram:byteenable2
	wire          mm_interconnect_2_ocram_s2_write;                                    // mm_interconnect_2:ocram_s2_write -> ocram:write2
	wire   [31:0] mm_interconnect_2_ocram_s2_writedata;                                // mm_interconnect_2:ocram_s2_writedata -> ocram:writedata2
	wire          mm_interconnect_2_ocram_s2_clken;                                    // mm_interconnect_2:ocram_s2_clken -> ocram:clken2
	wire   [31:0] jtag_hps_master_readdata;                                            // mm_interconnect_3:jtag_hps_master_readdata -> jtag_hps:master_readdata
	wire          jtag_hps_master_waitrequest;                                         // mm_interconnect_3:jtag_hps_master_waitrequest -> jtag_hps:master_waitrequest
	wire   [31:0] jtag_hps_master_address;                                             // jtag_hps:master_address -> mm_interconnect_3:jtag_hps_master_address
	wire          jtag_hps_master_read;                                                // jtag_hps:master_read -> mm_interconnect_3:jtag_hps_master_read
	wire    [3:0] jtag_hps_master_byteenable;                                          // jtag_hps:master_byteenable -> mm_interconnect_3:jtag_hps_master_byteenable
	wire          jtag_hps_master_readdatavalid;                                       // mm_interconnect_3:jtag_hps_master_readdatavalid -> jtag_hps:master_readdatavalid
	wire          jtag_hps_master_write;                                               // jtag_hps:master_write -> mm_interconnect_3:jtag_hps_master_write
	wire   [31:0] jtag_hps_master_writedata;                                           // jtag_hps:master_writedata -> mm_interconnect_3:jtag_hps_master_writedata
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awburst;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_awburst -> arm_hps:f2h_AWBURST
	wire    [4:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awuser;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_awuser -> arm_hps:f2h_AWUSER
	wire    [3:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arlen;                       // mm_interconnect_3:arm_hps_f2h_axi_slave_arlen -> arm_hps:f2h_ARLEN
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_wstrb;                       // mm_interconnect_3:arm_hps_f2h_axi_slave_wstrb -> arm_hps:f2h_WSTRB
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_wready;                      // arm_hps:f2h_WREADY -> mm_interconnect_3:arm_hps_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_rid;                         // arm_hps:f2h_RID -> mm_interconnect_3:arm_hps_f2h_axi_slave_rid
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_rready;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_rready -> arm_hps:f2h_RREADY
	wire    [3:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awlen;                       // mm_interconnect_3:arm_hps_f2h_axi_slave_awlen -> arm_hps:f2h_AWLEN
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_wid;                         // mm_interconnect_3:arm_hps_f2h_axi_slave_wid -> arm_hps:f2h_WID
	wire    [3:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arcache;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_arcache -> arm_hps:f2h_ARCACHE
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_wvalid;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_wvalid -> arm_hps:f2h_WVALID
	wire   [31:0] mm_interconnect_3_arm_hps_f2h_axi_slave_araddr;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_araddr -> arm_hps:f2h_ARADDR
	wire    [2:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arprot;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_arprot -> arm_hps:f2h_ARPROT
	wire    [2:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awprot;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_awprot -> arm_hps:f2h_AWPROT
	wire   [63:0] mm_interconnect_3_arm_hps_f2h_axi_slave_wdata;                       // mm_interconnect_3:arm_hps_f2h_axi_slave_wdata -> arm_hps:f2h_WDATA
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_arvalid;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_arvalid -> arm_hps:f2h_ARVALID
	wire    [3:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awcache;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_awcache -> arm_hps:f2h_AWCACHE
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arid;                        // mm_interconnect_3:arm_hps_f2h_axi_slave_arid -> arm_hps:f2h_ARID
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arlock;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_arlock -> arm_hps:f2h_ARLOCK
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awlock;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_awlock -> arm_hps:f2h_AWLOCK
	wire   [31:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awaddr;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_awaddr -> arm_hps:f2h_AWADDR
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_bresp;                       // arm_hps:f2h_BRESP -> mm_interconnect_3:arm_hps_f2h_axi_slave_bresp
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_arready;                     // arm_hps:f2h_ARREADY -> mm_interconnect_3:arm_hps_f2h_axi_slave_arready
	wire   [63:0] mm_interconnect_3_arm_hps_f2h_axi_slave_rdata;                       // arm_hps:f2h_RDATA -> mm_interconnect_3:arm_hps_f2h_axi_slave_rdata
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_awready;                     // arm_hps:f2h_AWREADY -> mm_interconnect_3:arm_hps_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arburst;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_arburst -> arm_hps:f2h_ARBURST
	wire    [2:0] mm_interconnect_3_arm_hps_f2h_axi_slave_arsize;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_arsize -> arm_hps:f2h_ARSIZE
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_bready;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_bready -> arm_hps:f2h_BREADY
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_rlast;                       // arm_hps:f2h_RLAST -> mm_interconnect_3:arm_hps_f2h_axi_slave_rlast
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_wlast;                       // mm_interconnect_3:arm_hps_f2h_axi_slave_wlast -> arm_hps:f2h_WLAST
	wire    [1:0] mm_interconnect_3_arm_hps_f2h_axi_slave_rresp;                       // arm_hps:f2h_RRESP -> mm_interconnect_3:arm_hps_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awid;                        // mm_interconnect_3:arm_hps_f2h_axi_slave_awid -> arm_hps:f2h_AWID
	wire    [7:0] mm_interconnect_3_arm_hps_f2h_axi_slave_bid;                         // arm_hps:f2h_BID -> mm_interconnect_3:arm_hps_f2h_axi_slave_bid
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_bvalid;                      // arm_hps:f2h_BVALID -> mm_interconnect_3:arm_hps_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_3_arm_hps_f2h_axi_slave_awsize;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_awsize -> arm_hps:f2h_AWSIZE
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_awvalid;                     // mm_interconnect_3:arm_hps_f2h_axi_slave_awvalid -> arm_hps:f2h_AWVALID
	wire    [4:0] mm_interconnect_3_arm_hps_f2h_axi_slave_aruser;                      // mm_interconnect_3:arm_hps_f2h_axi_slave_aruser -> arm_hps:f2h_ARUSER
	wire          mm_interconnect_3_arm_hps_f2h_axi_slave_rvalid;                      // arm_hps:f2h_RVALID -> mm_interconnect_3:arm_hps_f2h_axi_slave_rvalid
	wire          irq_mapper_receiver0_irq;                                            // IOPeripherals:buttons_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                            // AudioSubsystem:csr_irq_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                            // IOPeripherals:gpio0_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                            // IOPeripherals:gpio1_irq_irq -> irq_mapper:receiver3_irq
	wire          irq_mapper_receiver4_irq;                                            // IOPeripherals:irda_uart_irq_irq -> irq_mapper:receiver4_irq
	wire          irq_mapper_receiver5_irq;                                            // interval_timer:irq -> irq_mapper:receiver5_irq
	wire          irq_mapper_receiver6_irq;                                            // IOPeripherals:jtag_uart_irq_irq -> irq_mapper:receiver6_irq
	wire          irq_mapper_receiver7_irq;                                            // IOPeripherals:mandelbrot_irq_irq -> irq_mapper:receiver7_irq
	wire          irq_mapper_receiver8_irq;                                            // IOPeripherals:ps2_0_irq_irq -> irq_mapper:receiver8_irq
	wire          irq_mapper_receiver9_irq;                                            // IOPeripherals:ps2_1_irq_irq -> irq_mapper:receiver9_irq
	wire   [31:0] arm_hps_f2h_irq0_irq;                                                // irq_mapper:sender_irq -> arm_hps:f2h_irq_p0
	wire   [31:0] arm_hps_f2h_irq1_irq;                                                // irq_mapper_001:sender_irq -> arm_hps:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [AudioSubsystem:reset_reset_n, IOPeripherals:sys_reset_reset_n, baremetal:reset, interval_timer:reset_n, mm_interconnect_2:jtag_fpga_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:ocram_reset1_reset_bridge_in_reset_reset, mm_interconnect_3:jtag_hps_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:jtag_hps_master_translator_reset_reset_bridge_in_reset_reset, ocram:reset, rst_translator:in_reset, sdram:reset_n, sysid:reset_n]
	wire          rst_controller_reset_out_reset_req;                                  // rst_controller:reset_req -> [baremetal:reset_req, ocram:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> [mm_interconnect_2:arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_3:arm_hps_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]
	wire    [1:0] boot_from_fpga_value;                                                // port fragment

	Top_AudioSubsystem audiosubsystem (
		.audio_refclk_clk (audio_refclk_clk),                                // audio_refclk.clk
		.clk_clk          (system_ref_pll_outclk0_clk),                      //          clk.clk
		.csr_address      (mm_interconnect_2_audiosubsystem_csr_address),    //          csr.address
		.csr_readdata     (mm_interconnect_2_audiosubsystem_csr_readdata),   //             .readdata
		.csr_writedata    (mm_interconnect_2_audiosubsystem_csr_writedata),  //             .writedata
		.csr_write        (mm_interconnect_2_audiosubsystem_csr_write),      //             .write
		.csr_read         (mm_interconnect_2_audiosubsystem_csr_read),       //             .read
		.csr_byteenable   (mm_interconnect_2_audiosubsystem_csr_byteenable), //             .byteenable
		.csr_chipselect   (mm_interconnect_2_audiosubsystem_csr_chipselect), //             .chipselect
		.csr_irq_irq      (irq_mapper_receiver1_irq),                        //      csr_irq.irq
		.reset_reset_n    (~rst_controller_reset_out_reset),                 //        reset.reset_n
		.wm8731_bclk      (wm8731_bclk),                                     //       wm8731.bclk
		.wm8731_adclrck   (wm8731_adclrck),                                  //             .adclrck
		.wm8731_adcdat    (wm8731_adcdat),                                   //             .adcdat
		.wm8731_daclrck   (wm8731_daclrck),                                  //             .daclrck
		.wm8731_dacdat    (wm8731_dacdat),                                   //             .dacdat
		.wm8731_xck_clk   (wm8731_xck_clk)                                   //   wm8731_xck.clk
	);

	Top_IOPeripherals ioperipherals (
		.buttons_export               (buttons_export),                                               //        buttons.export
		.buttons_irq_irq              (irq_mapper_receiver0_irq),                                     //    buttons_irq.irq
		.ddr_read_read                (ioperipherals_ddr_read_read),                                  //       ddr_read.read
		.ddr_read_readdatavalid       (ioperipherals_ddr_read_readdatavalid),                         //               .readdatavalid
		.ddr_read_waitrequest         (ioperipherals_ddr_read_waitrequest),                           //               .waitrequest
		.ddr_read_readdata            (ioperipherals_ddr_read_readdata),                              //               .readdata
		.ddr_read_burstcount          (ioperipherals_ddr_read_burstcount),                            //               .burstcount
		.ddr_read_address             (ioperipherals_ddr_read_address),                               //               .address
		.ddr_write_write              (ioperipherals_ddr_write_write),                                //      ddr_write.write
		.ddr_write_waitrequest        (ioperipherals_ddr_write_waitrequest),                          //               .waitrequest
		.ddr_write_writedata          (ioperipherals_ddr_write_writedata),                            //               .writedata
		.ddr_write_byteenable         (ioperipherals_ddr_write_byteenable),                           //               .byteenable
		.ddr_write_burstcount         (ioperipherals_ddr_write_burstcount),                           //               .burstcount
		.ddr_write_address            (ioperipherals_ddr_write_address),                              //               .address
		.gpio0_export                 (gpio0_export),                                                 //          gpio0.export
		.gpio0_irq_irq                (irq_mapper_receiver2_irq),                                     //      gpio0_irq.irq
		.gpio1_export                 (gpio1_export),                                                 //          gpio1.export
		.gpio1_irq_irq                (irq_mapper_receiver3_irq),                                     //      gpio1_irq.irq
		.hex0_export                  (hex0_export),                                                  //           hex0.export
		.hex1_export                  (hex1_export),                                                  //           hex1.export
		.hex2_export                  (hex2_export),                                                  //           hex2.export
		.hex3_export                  (hex3_export),                                                  //           hex3.export
		.hex4_export                  (hex4_export),                                                  //           hex4.export
		.hex5_export                  (hex5_export),                                                  //           hex5.export
		.irda_uart_tx                 (irda_uart_tx),                                                 //      irda_uart.tx
		.irda_uart_rx                 (irda_uart_rx),                                                 //               .rx
		.irda_uart_irq_irq            (irq_mapper_receiver4_irq),                                     //  irda_uart_irq.irq
		.jtag_uart_irq_irq            (irq_mapper_receiver6_irq),                                     //  jtag_uart_irq.irq
		.leds_export                  (leds_export),                                                  //           leds.export
		.mandelbrot_irq_irq           (irq_mapper_receiver7_irq),                                     // mandelbrot_irq.irq
		.peripheral_map_waitrequest   (mm_interconnect_2_ioperipherals_peripheral_map_waitrequest),   // peripheral_map.waitrequest
		.peripheral_map_readdata      (mm_interconnect_2_ioperipherals_peripheral_map_readdata),      //               .readdata
		.peripheral_map_readdatavalid (mm_interconnect_2_ioperipherals_peripheral_map_readdatavalid), //               .readdatavalid
		.peripheral_map_burstcount    (mm_interconnect_2_ioperipherals_peripheral_map_burstcount),    //               .burstcount
		.peripheral_map_writedata     (mm_interconnect_2_ioperipherals_peripheral_map_writedata),     //               .writedata
		.peripheral_map_address       (mm_interconnect_2_ioperipherals_peripheral_map_address),       //               .address
		.peripheral_map_write         (mm_interconnect_2_ioperipherals_peripheral_map_write),         //               .write
		.peripheral_map_read          (mm_interconnect_2_ioperipherals_peripheral_map_read),          //               .read
		.peripheral_map_byteenable    (mm_interconnect_2_ioperipherals_peripheral_map_byteenable),    //               .byteenable
		.peripheral_map_debugaccess   (mm_interconnect_2_ioperipherals_peripheral_map_debugaccess),   //               .debugaccess
		.ps2_0_CLK                    (ps2_0_CLK),                                                    //          ps2_0.CLK
		.ps2_0_DAT                    (ps2_0_DAT),                                                    //               .DAT
		.ps2_0_irq_irq                (irq_mapper_receiver8_irq),                                     //      ps2_0_irq.irq
		.ps2_1_CLK                    (ps2_1_CLK),                                                    //          ps2_1.CLK
		.ps2_1_DAT                    (ps2_1_DAT),                                                    //               .DAT
		.ps2_1_irq_irq                (irq_mapper_receiver9_irq),                                     //      ps2_1_irq.irq
		.switches_export              (switches_export),                                              //       switches.export
		.sys_clk_clk                  (system_ref_pll_outclk0_clk),                                   //        sys_clk.clk
		.sys_reset_reset_n            (~rst_controller_reset_out_reset)                               //      sys_reset.reset_n
	);

	Top_VGASubsystem vgasubsystem (
		.char_buffer_control_slave_address    (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_address),    // char_buffer_control_slave.address
		.char_buffer_control_slave_byteenable (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_byteenable), //                          .byteenable
		.char_buffer_control_slave_chipselect (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_chipselect), //                          .chipselect
		.char_buffer_control_slave_read       (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_read),       //                          .read
		.char_buffer_control_slave_write      (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_write),      //                          .write
		.char_buffer_control_slave_writedata  (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_writedata),  //                          .writedata
		.char_buffer_control_slave_readdata   (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_readdata),   //                          .readdata
		.char_buffer_slave_byteenable         (mm_interconnect_2_vgasubsystem_char_buffer_slave_byteenable),         //         char_buffer_slave.byteenable
		.char_buffer_slave_chipselect         (mm_interconnect_2_vgasubsystem_char_buffer_slave_chipselect),         //                          .chipselect
		.char_buffer_slave_read               (mm_interconnect_2_vgasubsystem_char_buffer_slave_read),               //                          .read
		.char_buffer_slave_write              (mm_interconnect_2_vgasubsystem_char_buffer_slave_write),              //                          .write
		.char_buffer_slave_writedata          (mm_interconnect_2_vgasubsystem_char_buffer_slave_writedata),          //                          .writedata
		.char_buffer_slave_readdata           (mm_interconnect_2_vgasubsystem_char_buffer_slave_readdata),           //                          .readdata
		.char_buffer_slave_waitrequest        (mm_interconnect_2_vgasubsystem_char_buffer_slave_waitrequest),        //                          .waitrequest
		.char_buffer_slave_address            (mm_interconnect_2_vgasubsystem_char_buffer_slave_address),            //                          .address
		.pixel_dma_control_slave_address      (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_address),      //   pixel_dma_control_slave.address
		.pixel_dma_control_slave_byteenable   (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_byteenable),   //                          .byteenable
		.pixel_dma_control_slave_read         (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_read),         //                          .read
		.pixel_dma_control_slave_write        (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_write),        //                          .write
		.pixel_dma_control_slave_writedata    (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_writedata),    //                          .writedata
		.pixel_dma_control_slave_readdata     (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_readdata),     //                          .readdata
		.pixel_dma_master_readdatavalid       (vgasubsystem_pixel_dma_master_readdatavalid),                         //          pixel_dma_master.readdatavalid
		.pixel_dma_master_waitrequest         (vgasubsystem_pixel_dma_master_waitrequest),                           //                          .waitrequest
		.pixel_dma_master_address             (vgasubsystem_pixel_dma_master_address),                               //                          .address
		.pixel_dma_master_lock                (vgasubsystem_pixel_dma_master_lock),                                  //                          .lock
		.pixel_dma_master_read                (vgasubsystem_pixel_dma_master_read),                                  //                          .read
		.pixel_dma_master_readdata            (vgasubsystem_pixel_dma_master_readdata),                              //                          .readdata
		.sys_clk_clk                          (system_ref_pll_outclk0_clk),                                          //                   sys_clk.clk
		.sys_reset_reset_n                    (~system_reset_reset_out_reset),                                       //                 sys_reset.reset_n
		.vga_CLK                              (vga_CLK),                                                             //                       vga.CLK
		.vga_HS                               (vga_HS),                                                              //                          .HS
		.vga_VS                               (vga_VS),                                                              //                          .VS
		.vga_BLANK                            (vga_BLANK),                                                           //                          .BLANK
		.vga_SYNC                             (vga_SYNC),                                                            //                          .SYNC
		.vga_R                                (vga_R),                                                               //                          .R
		.vga_G                                (vga_G),                                                               //                          .G
		.vga_B                                (vga_B),                                                               //                          .B
		.vga_pll_ref_clk_clk                  (vga_refclk_clk),                                                      //           vga_pll_ref_clk.clk
		.vga_pll_ref_reset_reset              (system_reset_reset_out_reset)                                         //         vga_pll_ref_reset.reset
	);

	Top_arm_hps #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_hps (
		.f2h_boot_from_fpga_ready      (boot_from_fpga_constant_boot_from_fpga_ready),      // f2h_boot_from_fpga.boot_from_fpga_ready
		.f2h_boot_from_fpga_on_failure (boot_from_fpga_constant_boot_from_fpga_on_failure), //                   .boot_from_fpga_on_failure
		.mem_a                         (memory_mem_a),                                      //             memory.mem_a
		.mem_ba                        (memory_mem_ba),                                     //                   .mem_ba
		.mem_ck                        (memory_mem_ck),                                     //                   .mem_ck
		.mem_ck_n                      (memory_mem_ck_n),                                   //                   .mem_ck_n
		.mem_cke                       (memory_mem_cke),                                    //                   .mem_cke
		.mem_cs_n                      (memory_mem_cs_n),                                   //                   .mem_cs_n
		.mem_ras_n                     (memory_mem_ras_n),                                  //                   .mem_ras_n
		.mem_cas_n                     (memory_mem_cas_n),                                  //                   .mem_cas_n
		.mem_we_n                      (memory_mem_we_n),                                   //                   .mem_we_n
		.mem_reset_n                   (memory_mem_reset_n),                                //                   .mem_reset_n
		.mem_dq                        (memory_mem_dq),                                     //                   .mem_dq
		.mem_dqs                       (memory_mem_dqs),                                    //                   .mem_dqs
		.mem_dqs_n                     (memory_mem_dqs_n),                                  //                   .mem_dqs_n
		.mem_odt                       (memory_mem_odt),                                    //                   .mem_odt
		.mem_dm                        (memory_mem_dm),                                     //                   .mem_dm
		.oct_rzqin                     (memory_oct_rzqin),                                  //                   .oct_rzqin
		.hps_io_emac1_inst_TX_CLK      (hps_io_hps_io_emac1_inst_TX_CLK),                   //             hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0        (hps_io_hps_io_emac1_inst_TXD0),                     //                   .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1        (hps_io_hps_io_emac1_inst_TXD1),                     //                   .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2        (hps_io_hps_io_emac1_inst_TXD2),                     //                   .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3        (hps_io_hps_io_emac1_inst_TXD3),                     //                   .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0        (hps_io_hps_io_emac1_inst_RXD0),                     //                   .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO        (hps_io_hps_io_emac1_inst_MDIO),                     //                   .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC         (hps_io_hps_io_emac1_inst_MDC),                      //                   .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL      (hps_io_hps_io_emac1_inst_RX_CTL),                   //                   .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL      (hps_io_hps_io_emac1_inst_TX_CTL),                   //                   .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK      (hps_io_hps_io_emac1_inst_RX_CLK),                   //                   .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1        (hps_io_hps_io_emac1_inst_RXD1),                     //                   .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2        (hps_io_hps_io_emac1_inst_RXD2),                     //                   .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3        (hps_io_hps_io_emac1_inst_RXD3),                     //                   .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0          (hps_io_hps_io_qspi_inst_IO0),                       //                   .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1          (hps_io_hps_io_qspi_inst_IO1),                       //                   .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2          (hps_io_hps_io_qspi_inst_IO2),                       //                   .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3          (hps_io_hps_io_qspi_inst_IO3),                       //                   .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0          (hps_io_hps_io_qspi_inst_SS0),                       //                   .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK          (hps_io_hps_io_qspi_inst_CLK),                       //                   .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD          (hps_io_hps_io_sdio_inst_CMD),                       //                   .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0           (hps_io_hps_io_sdio_inst_D0),                        //                   .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1           (hps_io_hps_io_sdio_inst_D1),                        //                   .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK          (hps_io_hps_io_sdio_inst_CLK),                       //                   .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2           (hps_io_hps_io_sdio_inst_D2),                        //                   .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3           (hps_io_hps_io_sdio_inst_D3),                        //                   .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0           (hps_io_hps_io_usb1_inst_D0),                        //                   .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1           (hps_io_hps_io_usb1_inst_D1),                        //                   .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2           (hps_io_hps_io_usb1_inst_D2),                        //                   .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3           (hps_io_hps_io_usb1_inst_D3),                        //                   .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4           (hps_io_hps_io_usb1_inst_D4),                        //                   .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5           (hps_io_hps_io_usb1_inst_D5),                        //                   .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6           (hps_io_hps_io_usb1_inst_D6),                        //                   .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7           (hps_io_hps_io_usb1_inst_D7),                        //                   .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK          (hps_io_hps_io_usb1_inst_CLK),                       //                   .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP          (hps_io_hps_io_usb1_inst_STP),                       //                   .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR          (hps_io_hps_io_usb1_inst_DIR),                       //                   .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT          (hps_io_hps_io_usb1_inst_NXT),                       //                   .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK         (hps_io_hps_io_spim1_inst_CLK),                      //                   .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI        (hps_io_hps_io_spim1_inst_MOSI),                     //                   .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO        (hps_io_hps_io_spim1_inst_MISO),                     //                   .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0         (hps_io_hps_io_spim1_inst_SS0),                      //                   .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX          (hps_io_hps_io_uart0_inst_RX),                       //                   .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX          (hps_io_hps_io_uart0_inst_TX),                       //                   .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA          (hps_io_hps_io_i2c0_inst_SDA),                       //                   .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL          (hps_io_hps_io_i2c0_inst_SCL),                       //                   .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA          (hps_io_hps_io_i2c1_inst_SDA),                       //                   .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL          (hps_io_hps_io_i2c1_inst_SCL),                       //                   .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09       (hps_io_hps_io_gpio_inst_GPIO09),                    //                   .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35       (hps_io_hps_io_gpio_inst_GPIO35),                    //                   .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40       (hps_io_hps_io_gpio_inst_GPIO40),                    //                   .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41       (hps_io_hps_io_gpio_inst_GPIO41),                    //                   .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48       (hps_io_hps_io_gpio_inst_GPIO48),                    //                   .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53       (hps_io_hps_io_gpio_inst_GPIO53),                    //                   .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54       (hps_io_hps_io_gpio_inst_GPIO54),                    //                   .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61       (hps_io_hps_io_gpio_inst_GPIO61),                    //                   .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                     (arm_hps_h2f_reset_reset),                           //          h2f_reset.reset_n
		.f2h_sdram0_clk                (system_ref_pll_outclk0_clk),                        //   f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS            (ioperipherals_ddr_read_address),                    //    f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT         (ioperipherals_ddr_read_burstcount),                 //                   .burstcount
		.f2h_sdram0_WAITREQUEST        (ioperipherals_ddr_read_waitrequest),                //                   .waitrequest
		.f2h_sdram0_READDATA           (ioperipherals_ddr_read_readdata),                   //                   .readdata
		.f2h_sdram0_READDATAVALID      (ioperipherals_ddr_read_readdatavalid),              //                   .readdatavalid
		.f2h_sdram0_READ               (ioperipherals_ddr_read_read),                       //                   .read
		.f2h_sdram1_clk                (system_ref_pll_outclk0_clk),                        //   f2h_sdram1_clock.clk
		.f2h_sdram1_ADDRESS            (ioperipherals_ddr_write_address),                   //    f2h_sdram1_data.address
		.f2h_sdram1_BURSTCOUNT         (ioperipherals_ddr_write_burstcount),                //                   .burstcount
		.f2h_sdram1_WAITREQUEST        (ioperipherals_ddr_write_waitrequest),               //                   .waitrequest
		.f2h_sdram1_WRITEDATA          (ioperipherals_ddr_write_writedata),                 //                   .writedata
		.f2h_sdram1_BYTEENABLE         (ioperipherals_ddr_write_byteenable),                //                   .byteenable
		.f2h_sdram1_WRITE              (ioperipherals_ddr_write_write),                     //                   .write
		.h2f_axi_clk                   (system_ref_pll_outclk0_clk),                        //      h2f_axi_clock.clk
		.h2f_AWID                      (arm_hps_h2f_axi_master_awid),                       //     h2f_axi_master.awid
		.h2f_AWADDR                    (arm_hps_h2f_axi_master_awaddr),                     //                   .awaddr
		.h2f_AWLEN                     (arm_hps_h2f_axi_master_awlen),                      //                   .awlen
		.h2f_AWSIZE                    (arm_hps_h2f_axi_master_awsize),                     //                   .awsize
		.h2f_AWBURST                   (arm_hps_h2f_axi_master_awburst),                    //                   .awburst
		.h2f_AWLOCK                    (arm_hps_h2f_axi_master_awlock),                     //                   .awlock
		.h2f_AWCACHE                   (arm_hps_h2f_axi_master_awcache),                    //                   .awcache
		.h2f_AWPROT                    (arm_hps_h2f_axi_master_awprot),                     //                   .awprot
		.h2f_AWVALID                   (arm_hps_h2f_axi_master_awvalid),                    //                   .awvalid
		.h2f_AWREADY                   (arm_hps_h2f_axi_master_awready),                    //                   .awready
		.h2f_WID                       (arm_hps_h2f_axi_master_wid),                        //                   .wid
		.h2f_WDATA                     (arm_hps_h2f_axi_master_wdata),                      //                   .wdata
		.h2f_WSTRB                     (arm_hps_h2f_axi_master_wstrb),                      //                   .wstrb
		.h2f_WLAST                     (arm_hps_h2f_axi_master_wlast),                      //                   .wlast
		.h2f_WVALID                    (arm_hps_h2f_axi_master_wvalid),                     //                   .wvalid
		.h2f_WREADY                    (arm_hps_h2f_axi_master_wready),                     //                   .wready
		.h2f_BID                       (arm_hps_h2f_axi_master_bid),                        //                   .bid
		.h2f_BRESP                     (arm_hps_h2f_axi_master_bresp),                      //                   .bresp
		.h2f_BVALID                    (arm_hps_h2f_axi_master_bvalid),                     //                   .bvalid
		.h2f_BREADY                    (arm_hps_h2f_axi_master_bready),                     //                   .bready
		.h2f_ARID                      (arm_hps_h2f_axi_master_arid),                       //                   .arid
		.h2f_ARADDR                    (arm_hps_h2f_axi_master_araddr),                     //                   .araddr
		.h2f_ARLEN                     (arm_hps_h2f_axi_master_arlen),                      //                   .arlen
		.h2f_ARSIZE                    (arm_hps_h2f_axi_master_arsize),                     //                   .arsize
		.h2f_ARBURST                   (arm_hps_h2f_axi_master_arburst),                    //                   .arburst
		.h2f_ARLOCK                    (arm_hps_h2f_axi_master_arlock),                     //                   .arlock
		.h2f_ARCACHE                   (arm_hps_h2f_axi_master_arcache),                    //                   .arcache
		.h2f_ARPROT                    (arm_hps_h2f_axi_master_arprot),                     //                   .arprot
		.h2f_ARVALID                   (arm_hps_h2f_axi_master_arvalid),                    //                   .arvalid
		.h2f_ARREADY                   (arm_hps_h2f_axi_master_arready),                    //                   .arready
		.h2f_RID                       (arm_hps_h2f_axi_master_rid),                        //                   .rid
		.h2f_RDATA                     (arm_hps_h2f_axi_master_rdata),                      //                   .rdata
		.h2f_RRESP                     (arm_hps_h2f_axi_master_rresp),                      //                   .rresp
		.h2f_RLAST                     (arm_hps_h2f_axi_master_rlast),                      //                   .rlast
		.h2f_RVALID                    (arm_hps_h2f_axi_master_rvalid),                     //                   .rvalid
		.h2f_RREADY                    (arm_hps_h2f_axi_master_rready),                     //                   .rready
		.f2h_axi_clk                   (system_ref_pll_outclk0_clk),                        //      f2h_axi_clock.clk
		.f2h_AWID                      (mm_interconnect_3_arm_hps_f2h_axi_slave_awid),      //      f2h_axi_slave.awid
		.f2h_AWADDR                    (mm_interconnect_3_arm_hps_f2h_axi_slave_awaddr),    //                   .awaddr
		.f2h_AWLEN                     (mm_interconnect_3_arm_hps_f2h_axi_slave_awlen),     //                   .awlen
		.f2h_AWSIZE                    (mm_interconnect_3_arm_hps_f2h_axi_slave_awsize),    //                   .awsize
		.f2h_AWBURST                   (mm_interconnect_3_arm_hps_f2h_axi_slave_awburst),   //                   .awburst
		.f2h_AWLOCK                    (mm_interconnect_3_arm_hps_f2h_axi_slave_awlock),    //                   .awlock
		.f2h_AWCACHE                   (mm_interconnect_3_arm_hps_f2h_axi_slave_awcache),   //                   .awcache
		.f2h_AWPROT                    (mm_interconnect_3_arm_hps_f2h_axi_slave_awprot),    //                   .awprot
		.f2h_AWVALID                   (mm_interconnect_3_arm_hps_f2h_axi_slave_awvalid),   //                   .awvalid
		.f2h_AWREADY                   (mm_interconnect_3_arm_hps_f2h_axi_slave_awready),   //                   .awready
		.f2h_AWUSER                    (mm_interconnect_3_arm_hps_f2h_axi_slave_awuser),    //                   .awuser
		.f2h_WID                       (mm_interconnect_3_arm_hps_f2h_axi_slave_wid),       //                   .wid
		.f2h_WDATA                     (mm_interconnect_3_arm_hps_f2h_axi_slave_wdata),     //                   .wdata
		.f2h_WSTRB                     (mm_interconnect_3_arm_hps_f2h_axi_slave_wstrb),     //                   .wstrb
		.f2h_WLAST                     (mm_interconnect_3_arm_hps_f2h_axi_slave_wlast),     //                   .wlast
		.f2h_WVALID                    (mm_interconnect_3_arm_hps_f2h_axi_slave_wvalid),    //                   .wvalid
		.f2h_WREADY                    (mm_interconnect_3_arm_hps_f2h_axi_slave_wready),    //                   .wready
		.f2h_BID                       (mm_interconnect_3_arm_hps_f2h_axi_slave_bid),       //                   .bid
		.f2h_BRESP                     (mm_interconnect_3_arm_hps_f2h_axi_slave_bresp),     //                   .bresp
		.f2h_BVALID                    (mm_interconnect_3_arm_hps_f2h_axi_slave_bvalid),    //                   .bvalid
		.f2h_BREADY                    (mm_interconnect_3_arm_hps_f2h_axi_slave_bready),    //                   .bready
		.f2h_ARID                      (mm_interconnect_3_arm_hps_f2h_axi_slave_arid),      //                   .arid
		.f2h_ARADDR                    (mm_interconnect_3_arm_hps_f2h_axi_slave_araddr),    //                   .araddr
		.f2h_ARLEN                     (mm_interconnect_3_arm_hps_f2h_axi_slave_arlen),     //                   .arlen
		.f2h_ARSIZE                    (mm_interconnect_3_arm_hps_f2h_axi_slave_arsize),    //                   .arsize
		.f2h_ARBURST                   (mm_interconnect_3_arm_hps_f2h_axi_slave_arburst),   //                   .arburst
		.f2h_ARLOCK                    (mm_interconnect_3_arm_hps_f2h_axi_slave_arlock),    //                   .arlock
		.f2h_ARCACHE                   (mm_interconnect_3_arm_hps_f2h_axi_slave_arcache),   //                   .arcache
		.f2h_ARPROT                    (mm_interconnect_3_arm_hps_f2h_axi_slave_arprot),    //                   .arprot
		.f2h_ARVALID                   (mm_interconnect_3_arm_hps_f2h_axi_slave_arvalid),   //                   .arvalid
		.f2h_ARREADY                   (mm_interconnect_3_arm_hps_f2h_axi_slave_arready),   //                   .arready
		.f2h_ARUSER                    (mm_interconnect_3_arm_hps_f2h_axi_slave_aruser),    //                   .aruser
		.f2h_RID                       (mm_interconnect_3_arm_hps_f2h_axi_slave_rid),       //                   .rid
		.f2h_RDATA                     (mm_interconnect_3_arm_hps_f2h_axi_slave_rdata),     //                   .rdata
		.f2h_RRESP                     (mm_interconnect_3_arm_hps_f2h_axi_slave_rresp),     //                   .rresp
		.f2h_RLAST                     (mm_interconnect_3_arm_hps_f2h_axi_slave_rlast),     //                   .rlast
		.f2h_RVALID                    (mm_interconnect_3_arm_hps_f2h_axi_slave_rvalid),    //                   .rvalid
		.f2h_RREADY                    (mm_interconnect_3_arm_hps_f2h_axi_slave_rready),    //                   .rready
		.h2f_lw_axi_clk                (system_ref_pll_outclk0_clk),                        //   h2f_lw_axi_clock.clk
		.h2f_lw_AWID                   (arm_hps_h2f_lw_axi_master_awid),                    //  h2f_lw_axi_master.awid
		.h2f_lw_AWADDR                 (arm_hps_h2f_lw_axi_master_awaddr),                  //                   .awaddr
		.h2f_lw_AWLEN                  (arm_hps_h2f_lw_axi_master_awlen),                   //                   .awlen
		.h2f_lw_AWSIZE                 (arm_hps_h2f_lw_axi_master_awsize),                  //                   .awsize
		.h2f_lw_AWBURST                (arm_hps_h2f_lw_axi_master_awburst),                 //                   .awburst
		.h2f_lw_AWLOCK                 (arm_hps_h2f_lw_axi_master_awlock),                  //                   .awlock
		.h2f_lw_AWCACHE                (arm_hps_h2f_lw_axi_master_awcache),                 //                   .awcache
		.h2f_lw_AWPROT                 (arm_hps_h2f_lw_axi_master_awprot),                  //                   .awprot
		.h2f_lw_AWVALID                (arm_hps_h2f_lw_axi_master_awvalid),                 //                   .awvalid
		.h2f_lw_AWREADY                (arm_hps_h2f_lw_axi_master_awready),                 //                   .awready
		.h2f_lw_WID                    (arm_hps_h2f_lw_axi_master_wid),                     //                   .wid
		.h2f_lw_WDATA                  (arm_hps_h2f_lw_axi_master_wdata),                   //                   .wdata
		.h2f_lw_WSTRB                  (arm_hps_h2f_lw_axi_master_wstrb),                   //                   .wstrb
		.h2f_lw_WLAST                  (arm_hps_h2f_lw_axi_master_wlast),                   //                   .wlast
		.h2f_lw_WVALID                 (arm_hps_h2f_lw_axi_master_wvalid),                  //                   .wvalid
		.h2f_lw_WREADY                 (arm_hps_h2f_lw_axi_master_wready),                  //                   .wready
		.h2f_lw_BID                    (arm_hps_h2f_lw_axi_master_bid),                     //                   .bid
		.h2f_lw_BRESP                  (arm_hps_h2f_lw_axi_master_bresp),                   //                   .bresp
		.h2f_lw_BVALID                 (arm_hps_h2f_lw_axi_master_bvalid),                  //                   .bvalid
		.h2f_lw_BREADY                 (arm_hps_h2f_lw_axi_master_bready),                  //                   .bready
		.h2f_lw_ARID                   (arm_hps_h2f_lw_axi_master_arid),                    //                   .arid
		.h2f_lw_ARADDR                 (arm_hps_h2f_lw_axi_master_araddr),                  //                   .araddr
		.h2f_lw_ARLEN                  (arm_hps_h2f_lw_axi_master_arlen),                   //                   .arlen
		.h2f_lw_ARSIZE                 (arm_hps_h2f_lw_axi_master_arsize),                  //                   .arsize
		.h2f_lw_ARBURST                (arm_hps_h2f_lw_axi_master_arburst),                 //                   .arburst
		.h2f_lw_ARLOCK                 (arm_hps_h2f_lw_axi_master_arlock),                  //                   .arlock
		.h2f_lw_ARCACHE                (arm_hps_h2f_lw_axi_master_arcache),                 //                   .arcache
		.h2f_lw_ARPROT                 (arm_hps_h2f_lw_axi_master_arprot),                  //                   .arprot
		.h2f_lw_ARVALID                (arm_hps_h2f_lw_axi_master_arvalid),                 //                   .arvalid
		.h2f_lw_ARREADY                (arm_hps_h2f_lw_axi_master_arready),                 //                   .arready
		.h2f_lw_RID                    (arm_hps_h2f_lw_axi_master_rid),                     //                   .rid
		.h2f_lw_RDATA                  (arm_hps_h2f_lw_axi_master_rdata),                   //                   .rdata
		.h2f_lw_RRESP                  (arm_hps_h2f_lw_axi_master_rresp),                   //                   .rresp
		.h2f_lw_RLAST                  (arm_hps_h2f_lw_axi_master_rlast),                   //                   .rlast
		.h2f_lw_RVALID                 (arm_hps_h2f_lw_axi_master_rvalid),                  //                   .rvalid
		.h2f_lw_RREADY                 (arm_hps_h2f_lw_axi_master_rready),                  //                   .rready
		.f2h_irq_p0                    (arm_hps_f2h_irq0_irq),                              //           f2h_irq0.irq
		.f2h_irq_p1                    (arm_hps_f2h_irq1_irq)                               //           f2h_irq1.irq
	);

	Top_baremetal baremetal (
		.clk        (system_ref_pll_outclk0_clk),                //   clk1.clk
		.address    (mm_interconnect_2_baremetal_s1_address),    //     s1.address
		.clken      (mm_interconnect_2_baremetal_s1_clken),      //       .clken
		.chipselect (mm_interconnect_2_baremetal_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_2_baremetal_s1_write),      //       .write
		.readdata   (mm_interconnect_2_baremetal_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_2_baremetal_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_2_baremetal_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze     (1'b0)                                       // (terminated)
	);

	constant_num_multi_hw #(
		.VALUE ("00"),
		.WIDTH (2)
	) boot_from_fpga (
		.value ({boot_from_fpga_value[1],boot_from_fpga_value[0]})  // constant.boot_from_fpga_on_failure
	);

	Top_interval_timer interval_timer (
		.clk        (system_ref_pll_outclk0_clk),                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_2_interval_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_2_interval_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_2_interval_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_2_interval_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_2_interval_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                        //   irq.irq
	);

	Top_jtag_fpga #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_fpga (
		.clk_clk              (system_ref_pll_outclk0_clk),     //          clk.clk
		.clk_reset_reset      (system_reset_reset_out_reset),   //    clk_reset.reset
		.master_address       (jtag_fpga_master_address),       //       master.address
		.master_readdata      (jtag_fpga_master_readdata),      //             .readdata
		.master_read          (jtag_fpga_master_read),          //             .read
		.master_write         (jtag_fpga_master_write),         //             .write
		.master_writedata     (jtag_fpga_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_fpga_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_fpga_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_fpga_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                // master_reset.reset
	);

	Top_jtag_fpga #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) jtag_hps (
		.clk_clk              (system_ref_pll_outclk0_clk),    //          clk.clk
		.clk_reset_reset      (system_reset_reset_out_reset),  //    clk_reset.reset
		.master_address       (jtag_hps_master_address),       //       master.address
		.master_readdata      (jtag_hps_master_readdata),      //             .readdata
		.master_read          (jtag_hps_master_read),          //             .read
		.master_write         (jtag_hps_master_write),         //             .write
		.master_writedata     (jtag_hps_master_writedata),     //             .writedata
		.master_waitrequest   (jtag_hps_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (jtag_hps_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (jtag_hps_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	Top_ocram ocram (
		.address     (mm_interconnect_2_ocram_s1_address),    //     s1.address
		.clken       (mm_interconnect_2_ocram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_2_ocram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_2_ocram_s1_write),      //       .write
		.readdata    (mm_interconnect_2_ocram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_2_ocram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_2_ocram_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_2_ocram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_2_ocram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_2_ocram_s2_clken),      //       .clken
		.write2      (mm_interconnect_2_ocram_s2_write),      //       .write
		.readdata2   (mm_interconnect_2_ocram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_2_ocram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_2_ocram_s2_byteenable), //       .byteenable
		.clk         (system_ref_pll_outclk0_clk),            //   clk1.clk
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	pll_locked_to_reset_hw pll_locked (
		.locked  (system_ref_pll_locked_export), // locked.export
		.reset_n (pll_locked_reset_reset)        //  reset.reset_n
	);

	Top_sdram sdram (
		.clk            (system_ref_pll_outclk0_clk),               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_2_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_2_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_2_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_2_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_2_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_2_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_2_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_2_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_2_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	Top_sysid sysid (
		.clock    (system_ref_pll_outclk0_clk),                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_2_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_2_sysid_control_slave_address)   //              .address
	);

	Top_system_ref_pll system_ref_pll (
		.refclk   (system_ref_clk_clk),           //  refclk.clk
		.rst      (system_ref_reset_reset),       //   reset.reset
		.outclk_0 (system_ref_pll_outclk0_clk),   // outclk0.clk
		.outclk_1 (sdram_clk_clk),                // outclk1.clk
		.locked   (system_ref_pll_locked_export)  //  locked.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) system_reset (
		.reset_in0      (~pll_locked_reset_reset),      // reset_in0.reset
		.reset_in1      (~arm_hps_h2f_reset_reset),     // reset_in1.reset
		.clk            (system_ref_pll_outclk0_clk),   //       clk.clk
		.reset_out      (system_reset_reset_out_reset), // reset_out.reset
		.reset_req      (),                             // (terminated)
		.reset_req_in0  (1'b0),                         // (terminated)
		.reset_req_in1  (1'b0),                         // (terminated)
		.reset_in2      (1'b0),                         // (terminated)
		.reset_req_in2  (1'b0),                         // (terminated)
		.reset_in3      (1'b0),                         // (terminated)
		.reset_req_in3  (1'b0),                         // (terminated)
		.reset_in4      (1'b0),                         // (terminated)
		.reset_req_in4  (1'b0),                         // (terminated)
		.reset_in5      (1'b0),                         // (terminated)
		.reset_req_in5  (1'b0),                         // (terminated)
		.reset_in6      (1'b0),                         // (terminated)
		.reset_req_in6  (1'b0),                         // (terminated)
		.reset_in7      (1'b0),                         // (terminated)
		.reset_req_in7  (1'b0),                         // (terminated)
		.reset_in8      (1'b0),                         // (terminated)
		.reset_req_in8  (1'b0),                         // (terminated)
		.reset_in9      (1'b0),                         // (terminated)
		.reset_req_in9  (1'b0),                         // (terminated)
		.reset_in10     (1'b0),                         // (terminated)
		.reset_req_in10 (1'b0),                         // (terminated)
		.reset_in11     (1'b0),                         // (terminated)
		.reset_req_in11 (1'b0),                         // (terminated)
		.reset_in12     (1'b0),                         // (terminated)
		.reset_req_in12 (1'b0),                         // (terminated)
		.reset_in13     (1'b0),                         // (terminated)
		.reset_req_in13 (1'b0),                         // (terminated)
		.reset_in14     (1'b0),                         // (terminated)
		.reset_req_in14 (1'b0),                         // (terminated)
		.reset_in15     (1'b0),                         // (terminated)
		.reset_req_in15 (1'b0)                          // (terminated)
	);

	Top_mm_interconnect_2 mm_interconnect_2 (
		.arm_hps_h2f_axi_master_awid                                        (arm_hps_h2f_axi_master_awid),                                         //                                       arm_hps_h2f_axi_master.awid
		.arm_hps_h2f_axi_master_awaddr                                      (arm_hps_h2f_axi_master_awaddr),                                       //                                                             .awaddr
		.arm_hps_h2f_axi_master_awlen                                       (arm_hps_h2f_axi_master_awlen),                                        //                                                             .awlen
		.arm_hps_h2f_axi_master_awsize                                      (arm_hps_h2f_axi_master_awsize),                                       //                                                             .awsize
		.arm_hps_h2f_axi_master_awburst                                     (arm_hps_h2f_axi_master_awburst),                                      //                                                             .awburst
		.arm_hps_h2f_axi_master_awlock                                      (arm_hps_h2f_axi_master_awlock),                                       //                                                             .awlock
		.arm_hps_h2f_axi_master_awcache                                     (arm_hps_h2f_axi_master_awcache),                                      //                                                             .awcache
		.arm_hps_h2f_axi_master_awprot                                      (arm_hps_h2f_axi_master_awprot),                                       //                                                             .awprot
		.arm_hps_h2f_axi_master_awvalid                                     (arm_hps_h2f_axi_master_awvalid),                                      //                                                             .awvalid
		.arm_hps_h2f_axi_master_awready                                     (arm_hps_h2f_axi_master_awready),                                      //                                                             .awready
		.arm_hps_h2f_axi_master_wid                                         (arm_hps_h2f_axi_master_wid),                                          //                                                             .wid
		.arm_hps_h2f_axi_master_wdata                                       (arm_hps_h2f_axi_master_wdata),                                        //                                                             .wdata
		.arm_hps_h2f_axi_master_wstrb                                       (arm_hps_h2f_axi_master_wstrb),                                        //                                                             .wstrb
		.arm_hps_h2f_axi_master_wlast                                       (arm_hps_h2f_axi_master_wlast),                                        //                                                             .wlast
		.arm_hps_h2f_axi_master_wvalid                                      (arm_hps_h2f_axi_master_wvalid),                                       //                                                             .wvalid
		.arm_hps_h2f_axi_master_wready                                      (arm_hps_h2f_axi_master_wready),                                       //                                                             .wready
		.arm_hps_h2f_axi_master_bid                                         (arm_hps_h2f_axi_master_bid),                                          //                                                             .bid
		.arm_hps_h2f_axi_master_bresp                                       (arm_hps_h2f_axi_master_bresp),                                        //                                                             .bresp
		.arm_hps_h2f_axi_master_bvalid                                      (arm_hps_h2f_axi_master_bvalid),                                       //                                                             .bvalid
		.arm_hps_h2f_axi_master_bready                                      (arm_hps_h2f_axi_master_bready),                                       //                                                             .bready
		.arm_hps_h2f_axi_master_arid                                        (arm_hps_h2f_axi_master_arid),                                         //                                                             .arid
		.arm_hps_h2f_axi_master_araddr                                      (arm_hps_h2f_axi_master_araddr),                                       //                                                             .araddr
		.arm_hps_h2f_axi_master_arlen                                       (arm_hps_h2f_axi_master_arlen),                                        //                                                             .arlen
		.arm_hps_h2f_axi_master_arsize                                      (arm_hps_h2f_axi_master_arsize),                                       //                                                             .arsize
		.arm_hps_h2f_axi_master_arburst                                     (arm_hps_h2f_axi_master_arburst),                                      //                                                             .arburst
		.arm_hps_h2f_axi_master_arlock                                      (arm_hps_h2f_axi_master_arlock),                                       //                                                             .arlock
		.arm_hps_h2f_axi_master_arcache                                     (arm_hps_h2f_axi_master_arcache),                                      //                                                             .arcache
		.arm_hps_h2f_axi_master_arprot                                      (arm_hps_h2f_axi_master_arprot),                                       //                                                             .arprot
		.arm_hps_h2f_axi_master_arvalid                                     (arm_hps_h2f_axi_master_arvalid),                                      //                                                             .arvalid
		.arm_hps_h2f_axi_master_arready                                     (arm_hps_h2f_axi_master_arready),                                      //                                                             .arready
		.arm_hps_h2f_axi_master_rid                                         (arm_hps_h2f_axi_master_rid),                                          //                                                             .rid
		.arm_hps_h2f_axi_master_rdata                                       (arm_hps_h2f_axi_master_rdata),                                        //                                                             .rdata
		.arm_hps_h2f_axi_master_rresp                                       (arm_hps_h2f_axi_master_rresp),                                        //                                                             .rresp
		.arm_hps_h2f_axi_master_rlast                                       (arm_hps_h2f_axi_master_rlast),                                        //                                                             .rlast
		.arm_hps_h2f_axi_master_rvalid                                      (arm_hps_h2f_axi_master_rvalid),                                       //                                                             .rvalid
		.arm_hps_h2f_axi_master_rready                                      (arm_hps_h2f_axi_master_rready),                                       //                                                             .rready
		.arm_hps_h2f_lw_axi_master_awid                                     (arm_hps_h2f_lw_axi_master_awid),                                      //                                    arm_hps_h2f_lw_axi_master.awid
		.arm_hps_h2f_lw_axi_master_awaddr                                   (arm_hps_h2f_lw_axi_master_awaddr),                                    //                                                             .awaddr
		.arm_hps_h2f_lw_axi_master_awlen                                    (arm_hps_h2f_lw_axi_master_awlen),                                     //                                                             .awlen
		.arm_hps_h2f_lw_axi_master_awsize                                   (arm_hps_h2f_lw_axi_master_awsize),                                    //                                                             .awsize
		.arm_hps_h2f_lw_axi_master_awburst                                  (arm_hps_h2f_lw_axi_master_awburst),                                   //                                                             .awburst
		.arm_hps_h2f_lw_axi_master_awlock                                   (arm_hps_h2f_lw_axi_master_awlock),                                    //                                                             .awlock
		.arm_hps_h2f_lw_axi_master_awcache                                  (arm_hps_h2f_lw_axi_master_awcache),                                   //                                                             .awcache
		.arm_hps_h2f_lw_axi_master_awprot                                   (arm_hps_h2f_lw_axi_master_awprot),                                    //                                                             .awprot
		.arm_hps_h2f_lw_axi_master_awvalid                                  (arm_hps_h2f_lw_axi_master_awvalid),                                   //                                                             .awvalid
		.arm_hps_h2f_lw_axi_master_awready                                  (arm_hps_h2f_lw_axi_master_awready),                                   //                                                             .awready
		.arm_hps_h2f_lw_axi_master_wid                                      (arm_hps_h2f_lw_axi_master_wid),                                       //                                                             .wid
		.arm_hps_h2f_lw_axi_master_wdata                                    (arm_hps_h2f_lw_axi_master_wdata),                                     //                                                             .wdata
		.arm_hps_h2f_lw_axi_master_wstrb                                    (arm_hps_h2f_lw_axi_master_wstrb),                                     //                                                             .wstrb
		.arm_hps_h2f_lw_axi_master_wlast                                    (arm_hps_h2f_lw_axi_master_wlast),                                     //                                                             .wlast
		.arm_hps_h2f_lw_axi_master_wvalid                                   (arm_hps_h2f_lw_axi_master_wvalid),                                    //                                                             .wvalid
		.arm_hps_h2f_lw_axi_master_wready                                   (arm_hps_h2f_lw_axi_master_wready),                                    //                                                             .wready
		.arm_hps_h2f_lw_axi_master_bid                                      (arm_hps_h2f_lw_axi_master_bid),                                       //                                                             .bid
		.arm_hps_h2f_lw_axi_master_bresp                                    (arm_hps_h2f_lw_axi_master_bresp),                                     //                                                             .bresp
		.arm_hps_h2f_lw_axi_master_bvalid                                   (arm_hps_h2f_lw_axi_master_bvalid),                                    //                                                             .bvalid
		.arm_hps_h2f_lw_axi_master_bready                                   (arm_hps_h2f_lw_axi_master_bready),                                    //                                                             .bready
		.arm_hps_h2f_lw_axi_master_arid                                     (arm_hps_h2f_lw_axi_master_arid),                                      //                                                             .arid
		.arm_hps_h2f_lw_axi_master_araddr                                   (arm_hps_h2f_lw_axi_master_araddr),                                    //                                                             .araddr
		.arm_hps_h2f_lw_axi_master_arlen                                    (arm_hps_h2f_lw_axi_master_arlen),                                     //                                                             .arlen
		.arm_hps_h2f_lw_axi_master_arsize                                   (arm_hps_h2f_lw_axi_master_arsize),                                    //                                                             .arsize
		.arm_hps_h2f_lw_axi_master_arburst                                  (arm_hps_h2f_lw_axi_master_arburst),                                   //                                                             .arburst
		.arm_hps_h2f_lw_axi_master_arlock                                   (arm_hps_h2f_lw_axi_master_arlock),                                    //                                                             .arlock
		.arm_hps_h2f_lw_axi_master_arcache                                  (arm_hps_h2f_lw_axi_master_arcache),                                   //                                                             .arcache
		.arm_hps_h2f_lw_axi_master_arprot                                   (arm_hps_h2f_lw_axi_master_arprot),                                    //                                                             .arprot
		.arm_hps_h2f_lw_axi_master_arvalid                                  (arm_hps_h2f_lw_axi_master_arvalid),                                   //                                                             .arvalid
		.arm_hps_h2f_lw_axi_master_arready                                  (arm_hps_h2f_lw_axi_master_arready),                                   //                                                             .arready
		.arm_hps_h2f_lw_axi_master_rid                                      (arm_hps_h2f_lw_axi_master_rid),                                       //                                                             .rid
		.arm_hps_h2f_lw_axi_master_rdata                                    (arm_hps_h2f_lw_axi_master_rdata),                                     //                                                             .rdata
		.arm_hps_h2f_lw_axi_master_rresp                                    (arm_hps_h2f_lw_axi_master_rresp),                                     //                                                             .rresp
		.arm_hps_h2f_lw_axi_master_rlast                                    (arm_hps_h2f_lw_axi_master_rlast),                                     //                                                             .rlast
		.arm_hps_h2f_lw_axi_master_rvalid                                   (arm_hps_h2f_lw_axi_master_rvalid),                                    //                                                             .rvalid
		.arm_hps_h2f_lw_axi_master_rready                                   (arm_hps_h2f_lw_axi_master_rready),                                    //                                                             .rready
		.system_ref_pll_outclk0_clk                                         (system_ref_pll_outclk0_clk),                                          //                                       system_ref_pll_outclk0.clk
		.arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                                  // arm_hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.jtag_fpga_clk_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                                      //                    jtag_fpga_clk_reset_reset_bridge_in_reset.reset
		.ocram_reset1_reset_bridge_in_reset_reset                           (rst_controller_reset_out_reset),                                      //                           ocram_reset1_reset_bridge_in_reset.reset
		.jtag_fpga_master_address                                           (jtag_fpga_master_address),                                            //                                             jtag_fpga_master.address
		.jtag_fpga_master_waitrequest                                       (jtag_fpga_master_waitrequest),                                        //                                                             .waitrequest
		.jtag_fpga_master_byteenable                                        (jtag_fpga_master_byteenable),                                         //                                                             .byteenable
		.jtag_fpga_master_read                                              (jtag_fpga_master_read),                                               //                                                             .read
		.jtag_fpga_master_readdata                                          (jtag_fpga_master_readdata),                                           //                                                             .readdata
		.jtag_fpga_master_readdatavalid                                     (jtag_fpga_master_readdatavalid),                                      //                                                             .readdatavalid
		.jtag_fpga_master_write                                             (jtag_fpga_master_write),                                              //                                                             .write
		.jtag_fpga_master_writedata                                         (jtag_fpga_master_writedata),                                          //                                                             .writedata
		.VGASubsystem_pixel_dma_master_address                              (vgasubsystem_pixel_dma_master_address),                               //                                VGASubsystem_pixel_dma_master.address
		.VGASubsystem_pixel_dma_master_waitrequest                          (vgasubsystem_pixel_dma_master_waitrequest),                           //                                                             .waitrequest
		.VGASubsystem_pixel_dma_master_read                                 (vgasubsystem_pixel_dma_master_read),                                  //                                                             .read
		.VGASubsystem_pixel_dma_master_readdata                             (vgasubsystem_pixel_dma_master_readdata),                              //                                                             .readdata
		.VGASubsystem_pixel_dma_master_readdatavalid                        (vgasubsystem_pixel_dma_master_readdatavalid),                         //                                                             .readdatavalid
		.VGASubsystem_pixel_dma_master_lock                                 (vgasubsystem_pixel_dma_master_lock),                                  //                                                             .lock
		.AudioSubsystem_csr_address                                         (mm_interconnect_2_audiosubsystem_csr_address),                        //                                           AudioSubsystem_csr.address
		.AudioSubsystem_csr_write                                           (mm_interconnect_2_audiosubsystem_csr_write),                          //                                                             .write
		.AudioSubsystem_csr_read                                            (mm_interconnect_2_audiosubsystem_csr_read),                           //                                                             .read
		.AudioSubsystem_csr_readdata                                        (mm_interconnect_2_audiosubsystem_csr_readdata),                       //                                                             .readdata
		.AudioSubsystem_csr_writedata                                       (mm_interconnect_2_audiosubsystem_csr_writedata),                      //                                                             .writedata
		.AudioSubsystem_csr_byteenable                                      (mm_interconnect_2_audiosubsystem_csr_byteenable),                     //                                                             .byteenable
		.AudioSubsystem_csr_chipselect                                      (mm_interconnect_2_audiosubsystem_csr_chipselect),                     //                                                             .chipselect
		.baremetal_s1_address                                               (mm_interconnect_2_baremetal_s1_address),                              //                                                 baremetal_s1.address
		.baremetal_s1_write                                                 (mm_interconnect_2_baremetal_s1_write),                                //                                                             .write
		.baremetal_s1_readdata                                              (mm_interconnect_2_baremetal_s1_readdata),                             //                                                             .readdata
		.baremetal_s1_writedata                                             (mm_interconnect_2_baremetal_s1_writedata),                            //                                                             .writedata
		.baremetal_s1_byteenable                                            (mm_interconnect_2_baremetal_s1_byteenable),                           //                                                             .byteenable
		.baremetal_s1_chipselect                                            (mm_interconnect_2_baremetal_s1_chipselect),                           //                                                             .chipselect
		.baremetal_s1_clken                                                 (mm_interconnect_2_baremetal_s1_clken),                                //                                                             .clken
		.interval_timer_s1_address                                          (mm_interconnect_2_interval_timer_s1_address),                         //                                            interval_timer_s1.address
		.interval_timer_s1_write                                            (mm_interconnect_2_interval_timer_s1_write),                           //                                                             .write
		.interval_timer_s1_readdata                                         (mm_interconnect_2_interval_timer_s1_readdata),                        //                                                             .readdata
		.interval_timer_s1_writedata                                        (mm_interconnect_2_interval_timer_s1_writedata),                       //                                                             .writedata
		.interval_timer_s1_chipselect                                       (mm_interconnect_2_interval_timer_s1_chipselect),                      //                                                             .chipselect
		.IOPeripherals_peripheral_map_address                               (mm_interconnect_2_ioperipherals_peripheral_map_address),              //                                 IOPeripherals_peripheral_map.address
		.IOPeripherals_peripheral_map_write                                 (mm_interconnect_2_ioperipherals_peripheral_map_write),                //                                                             .write
		.IOPeripherals_peripheral_map_read                                  (mm_interconnect_2_ioperipherals_peripheral_map_read),                 //                                                             .read
		.IOPeripherals_peripheral_map_readdata                              (mm_interconnect_2_ioperipherals_peripheral_map_readdata),             //                                                             .readdata
		.IOPeripherals_peripheral_map_writedata                             (mm_interconnect_2_ioperipherals_peripheral_map_writedata),            //                                                             .writedata
		.IOPeripherals_peripheral_map_burstcount                            (mm_interconnect_2_ioperipherals_peripheral_map_burstcount),           //                                                             .burstcount
		.IOPeripherals_peripheral_map_byteenable                            (mm_interconnect_2_ioperipherals_peripheral_map_byteenable),           //                                                             .byteenable
		.IOPeripherals_peripheral_map_readdatavalid                         (mm_interconnect_2_ioperipherals_peripheral_map_readdatavalid),        //                                                             .readdatavalid
		.IOPeripherals_peripheral_map_waitrequest                           (mm_interconnect_2_ioperipherals_peripheral_map_waitrequest),          //                                                             .waitrequest
		.IOPeripherals_peripheral_map_debugaccess                           (mm_interconnect_2_ioperipherals_peripheral_map_debugaccess),          //                                                             .debugaccess
		.ocram_s1_address                                                   (mm_interconnect_2_ocram_s1_address),                                  //                                                     ocram_s1.address
		.ocram_s1_write                                                     (mm_interconnect_2_ocram_s1_write),                                    //                                                             .write
		.ocram_s1_readdata                                                  (mm_interconnect_2_ocram_s1_readdata),                                 //                                                             .readdata
		.ocram_s1_writedata                                                 (mm_interconnect_2_ocram_s1_writedata),                                //                                                             .writedata
		.ocram_s1_byteenable                                                (mm_interconnect_2_ocram_s1_byteenable),                               //                                                             .byteenable
		.ocram_s1_chipselect                                                (mm_interconnect_2_ocram_s1_chipselect),                               //                                                             .chipselect
		.ocram_s1_clken                                                     (mm_interconnect_2_ocram_s1_clken),                                    //                                                             .clken
		.ocram_s2_address                                                   (mm_interconnect_2_ocram_s2_address),                                  //                                                     ocram_s2.address
		.ocram_s2_write                                                     (mm_interconnect_2_ocram_s2_write),                                    //                                                             .write
		.ocram_s2_readdata                                                  (mm_interconnect_2_ocram_s2_readdata),                                 //                                                             .readdata
		.ocram_s2_writedata                                                 (mm_interconnect_2_ocram_s2_writedata),                                //                                                             .writedata
		.ocram_s2_byteenable                                                (mm_interconnect_2_ocram_s2_byteenable),                               //                                                             .byteenable
		.ocram_s2_chipselect                                                (mm_interconnect_2_ocram_s2_chipselect),                               //                                                             .chipselect
		.ocram_s2_clken                                                     (mm_interconnect_2_ocram_s2_clken),                                    //                                                             .clken
		.sdram_s1_address                                                   (mm_interconnect_2_sdram_s1_address),                                  //                                                     sdram_s1.address
		.sdram_s1_write                                                     (mm_interconnect_2_sdram_s1_write),                                    //                                                             .write
		.sdram_s1_read                                                      (mm_interconnect_2_sdram_s1_read),                                     //                                                             .read
		.sdram_s1_readdata                                                  (mm_interconnect_2_sdram_s1_readdata),                                 //                                                             .readdata
		.sdram_s1_writedata                                                 (mm_interconnect_2_sdram_s1_writedata),                                //                                                             .writedata
		.sdram_s1_byteenable                                                (mm_interconnect_2_sdram_s1_byteenable),                               //                                                             .byteenable
		.sdram_s1_readdatavalid                                             (mm_interconnect_2_sdram_s1_readdatavalid),                            //                                                             .readdatavalid
		.sdram_s1_waitrequest                                               (mm_interconnect_2_sdram_s1_waitrequest),                              //                                                             .waitrequest
		.sdram_s1_chipselect                                                (mm_interconnect_2_sdram_s1_chipselect),                               //                                                             .chipselect
		.sysid_control_slave_address                                        (mm_interconnect_2_sysid_control_slave_address),                       //                                          sysid_control_slave.address
		.sysid_control_slave_readdata                                       (mm_interconnect_2_sysid_control_slave_readdata),                      //                                                             .readdata
		.VGASubsystem_char_buffer_control_slave_address                     (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_address),    //                       VGASubsystem_char_buffer_control_slave.address
		.VGASubsystem_char_buffer_control_slave_write                       (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_write),      //                                                             .write
		.VGASubsystem_char_buffer_control_slave_read                        (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_read),       //                                                             .read
		.VGASubsystem_char_buffer_control_slave_readdata                    (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_readdata),   //                                                             .readdata
		.VGASubsystem_char_buffer_control_slave_writedata                   (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_writedata),  //                                                             .writedata
		.VGASubsystem_char_buffer_control_slave_byteenable                  (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_byteenable), //                                                             .byteenable
		.VGASubsystem_char_buffer_control_slave_chipselect                  (mm_interconnect_2_vgasubsystem_char_buffer_control_slave_chipselect), //                                                             .chipselect
		.VGASubsystem_char_buffer_slave_address                             (mm_interconnect_2_vgasubsystem_char_buffer_slave_address),            //                               VGASubsystem_char_buffer_slave.address
		.VGASubsystem_char_buffer_slave_write                               (mm_interconnect_2_vgasubsystem_char_buffer_slave_write),              //                                                             .write
		.VGASubsystem_char_buffer_slave_read                                (mm_interconnect_2_vgasubsystem_char_buffer_slave_read),               //                                                             .read
		.VGASubsystem_char_buffer_slave_readdata                            (mm_interconnect_2_vgasubsystem_char_buffer_slave_readdata),           //                                                             .readdata
		.VGASubsystem_char_buffer_slave_writedata                           (mm_interconnect_2_vgasubsystem_char_buffer_slave_writedata),          //                                                             .writedata
		.VGASubsystem_char_buffer_slave_byteenable                          (mm_interconnect_2_vgasubsystem_char_buffer_slave_byteenable),         //                                                             .byteenable
		.VGASubsystem_char_buffer_slave_waitrequest                         (mm_interconnect_2_vgasubsystem_char_buffer_slave_waitrequest),        //                                                             .waitrequest
		.VGASubsystem_char_buffer_slave_chipselect                          (mm_interconnect_2_vgasubsystem_char_buffer_slave_chipselect),         //                                                             .chipselect
		.VGASubsystem_pixel_dma_control_slave_address                       (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_address),      //                         VGASubsystem_pixel_dma_control_slave.address
		.VGASubsystem_pixel_dma_control_slave_write                         (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_write),        //                                                             .write
		.VGASubsystem_pixel_dma_control_slave_read                          (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_read),         //                                                             .read
		.VGASubsystem_pixel_dma_control_slave_readdata                      (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_readdata),     //                                                             .readdata
		.VGASubsystem_pixel_dma_control_slave_writedata                     (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_writedata),    //                                                             .writedata
		.VGASubsystem_pixel_dma_control_slave_byteenable                    (mm_interconnect_2_vgasubsystem_pixel_dma_control_slave_byteenable)    //                                                             .byteenable
	);

	Top_mm_interconnect_3 mm_interconnect_3 (
		.arm_hps_f2h_axi_slave_awid                                         (mm_interconnect_3_arm_hps_f2h_axi_slave_awid),    //                                        arm_hps_f2h_axi_slave.awid
		.arm_hps_f2h_axi_slave_awaddr                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_awaddr),  //                                                             .awaddr
		.arm_hps_f2h_axi_slave_awlen                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_awlen),   //                                                             .awlen
		.arm_hps_f2h_axi_slave_awsize                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_awsize),  //                                                             .awsize
		.arm_hps_f2h_axi_slave_awburst                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_awburst), //                                                             .awburst
		.arm_hps_f2h_axi_slave_awlock                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_awlock),  //                                                             .awlock
		.arm_hps_f2h_axi_slave_awcache                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_awcache), //                                                             .awcache
		.arm_hps_f2h_axi_slave_awprot                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_awprot),  //                                                             .awprot
		.arm_hps_f2h_axi_slave_awuser                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_awuser),  //                                                             .awuser
		.arm_hps_f2h_axi_slave_awvalid                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_awvalid), //                                                             .awvalid
		.arm_hps_f2h_axi_slave_awready                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_awready), //                                                             .awready
		.arm_hps_f2h_axi_slave_wid                                          (mm_interconnect_3_arm_hps_f2h_axi_slave_wid),     //                                                             .wid
		.arm_hps_f2h_axi_slave_wdata                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_wdata),   //                                                             .wdata
		.arm_hps_f2h_axi_slave_wstrb                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_wstrb),   //                                                             .wstrb
		.arm_hps_f2h_axi_slave_wlast                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_wlast),   //                                                             .wlast
		.arm_hps_f2h_axi_slave_wvalid                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_wvalid),  //                                                             .wvalid
		.arm_hps_f2h_axi_slave_wready                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_wready),  //                                                             .wready
		.arm_hps_f2h_axi_slave_bid                                          (mm_interconnect_3_arm_hps_f2h_axi_slave_bid),     //                                                             .bid
		.arm_hps_f2h_axi_slave_bresp                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_bresp),   //                                                             .bresp
		.arm_hps_f2h_axi_slave_bvalid                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_bvalid),  //                                                             .bvalid
		.arm_hps_f2h_axi_slave_bready                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_bready),  //                                                             .bready
		.arm_hps_f2h_axi_slave_arid                                         (mm_interconnect_3_arm_hps_f2h_axi_slave_arid),    //                                                             .arid
		.arm_hps_f2h_axi_slave_araddr                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_araddr),  //                                                             .araddr
		.arm_hps_f2h_axi_slave_arlen                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_arlen),   //                                                             .arlen
		.arm_hps_f2h_axi_slave_arsize                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_arsize),  //                                                             .arsize
		.arm_hps_f2h_axi_slave_arburst                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_arburst), //                                                             .arburst
		.arm_hps_f2h_axi_slave_arlock                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_arlock),  //                                                             .arlock
		.arm_hps_f2h_axi_slave_arcache                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_arcache), //                                                             .arcache
		.arm_hps_f2h_axi_slave_arprot                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_arprot),  //                                                             .arprot
		.arm_hps_f2h_axi_slave_aruser                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_aruser),  //                                                             .aruser
		.arm_hps_f2h_axi_slave_arvalid                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_arvalid), //                                                             .arvalid
		.arm_hps_f2h_axi_slave_arready                                      (mm_interconnect_3_arm_hps_f2h_axi_slave_arready), //                                                             .arready
		.arm_hps_f2h_axi_slave_rid                                          (mm_interconnect_3_arm_hps_f2h_axi_slave_rid),     //                                                             .rid
		.arm_hps_f2h_axi_slave_rdata                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_rdata),   //                                                             .rdata
		.arm_hps_f2h_axi_slave_rresp                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_rresp),   //                                                             .rresp
		.arm_hps_f2h_axi_slave_rlast                                        (mm_interconnect_3_arm_hps_f2h_axi_slave_rlast),   //                                                             .rlast
		.arm_hps_f2h_axi_slave_rvalid                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_rvalid),  //                                                             .rvalid
		.arm_hps_f2h_axi_slave_rready                                       (mm_interconnect_3_arm_hps_f2h_axi_slave_rready),  //                                                             .rready
		.system_ref_pll_outclk0_clk                                         (system_ref_pll_outclk0_clk),                      //                                       system_ref_pll_outclk0.clk
		.arm_hps_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),              // arm_hps_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.jtag_hps_clk_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                  //                     jtag_hps_clk_reset_reset_bridge_in_reset.reset
		.jtag_hps_master_translator_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                  //       jtag_hps_master_translator_reset_reset_bridge_in_reset.reset
		.jtag_hps_master_address                                            (jtag_hps_master_address),                         //                                              jtag_hps_master.address
		.jtag_hps_master_waitrequest                                        (jtag_hps_master_waitrequest),                     //                                                             .waitrequest
		.jtag_hps_master_byteenable                                         (jtag_hps_master_byteenable),                      //                                                             .byteenable
		.jtag_hps_master_read                                               (jtag_hps_master_read),                            //                                                             .read
		.jtag_hps_master_readdata                                           (jtag_hps_master_readdata),                        //                                                             .readdata
		.jtag_hps_master_readdatavalid                                      (jtag_hps_master_readdatavalid),                   //                                                             .readdatavalid
		.jtag_hps_master_write                                              (jtag_hps_master_write),                           //                                                             .write
		.jtag_hps_master_writedata                                          (jtag_hps_master_writedata)                        //                                                             .writedata
	);

	Top_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq), // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq), // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq), // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq), // receiver9.irq
		.sender_irq    (arm_hps_f2h_irq0_irq)      //    sender.irq
	);

	Top_irq_mapper_001 irq_mapper_001 (
		.clk        (),                     //       clk.clk
		.reset      (),                     // clk_reset.reset
		.sender_irq (arm_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (system_reset_reset_out_reset),       // reset_in0.reset
		.clk            (system_ref_pll_outclk0_clk),         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (system_ref_pll_outclk0_clk),         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign boot_from_fpga_constant_boot_from_fpga_on_failure = { boot_from_fpga_value[0] };

	assign boot_from_fpga_constant_boot_from_fpga_ready = { boot_from_fpga_value[1] };

endmodule
